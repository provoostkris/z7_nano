

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-------------------------------------------------------------------------------
package ascii_pkg is

  -- create arrays for pixel map stores
  type t_xx08_arr  is array (natural range <>) of std_logic_vector(8-1 downto 0);     -- one row  in xx08 size
  type t_1608_arr  is array (natural range <>) of t_xx08_arr(0 to 15);                -- one char in 1608 size

  constant c_ascii_1608 : t_1608_arr( 0 to 94) :=
  (
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"), --! " ",0*/
  (x"00",x"00",x"00",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"00",x"00",x"18",x"18",x"00",x"00"), --! "!",1*/
  (x"00",x"48",x"6C",x"24",x"12",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"), --! """,2*/
  (x"00",x"00",x"00",x"24",x"24",x"24",x"7F",x"12",x"12",x"12",x"7F",x"12",x"12",x"12",x"00",x"00"), --! "#",3*/
  (x"00",x"00",x"08",x"1C",x"2A",x"2A",x"0A",x"0C",x"18",x"28",x"28",x"2A",x"2A",x"1C",x"08",x"08"), --! "$",4*/
  (x"00",x"00",x"00",x"22",x"25",x"15",x"15",x"15",x"2A",x"58",x"54",x"54",x"54",x"22",x"00",x"00"), --! "%",5*/
  (x"00",x"00",x"00",x"0C",x"12",x"12",x"12",x"0A",x"76",x"25",x"29",x"11",x"91",x"6E",x"00",x"00"), --! "&",6*/
  (x"00",x"06",x"06",x"04",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"), --! "'",7*/
  (x"00",x"40",x"20",x"10",x"10",x"08",x"08",x"08",x"08",x"08",x"08",x"10",x"10",x"20",x"40",x"00"), --! "(",8*/
  (x"00",x"02",x"04",x"08",x"08",x"10",x"10",x"10",x"10",x"10",x"10",x"08",x"08",x"04",x"02",x"00"), --! ")",9*/
  (x"00",x"00",x"00",x"00",x"08",x"08",x"6B",x"1C",x"1C",x"6B",x"08",x"08",x"00",x"00",x"00",x"00"), --! "*",10*/
  (x"00",x"00",x"00",x"00",x"08",x"08",x"08",x"08",x"7F",x"08",x"08",x"08",x"08",x"00",x"00",x"00"), --! "+",11*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"04",x"03"), --! ",",12*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00"), --! "-",13*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00"), --! ".",14*/
  (x"00",x"00",x"80",x"40",x"40",x"20",x"20",x"10",x"10",x"08",x"08",x"04",x"04",x"02",x"02",x"00"), --! "/",15*/
  (x"00",x"00",x"00",x"18",x"24",x"42",x"42",x"42",x"42",x"42",x"42",x"42",x"24",x"18",x"00",x"00"), --! "0",16*/
  (x"00",x"00",x"00",x"08",x"0E",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"3E",x"00",x"00"), --! "1",17*/
  (x"00",x"00",x"00",x"3C",x"42",x"42",x"42",x"20",x"20",x"10",x"08",x"04",x"42",x"7E",x"00",x"00"), --! "2",18*/
  (x"00",x"00",x"00",x"3C",x"42",x"42",x"20",x"18",x"20",x"40",x"40",x"42",x"22",x"1C",x"00",x"00"), --! "3",19*/
  (x"00",x"00",x"00",x"20",x"30",x"28",x"24",x"24",x"22",x"22",x"7E",x"20",x"20",x"78",x"00",x"00"), --! "4",20*/
  (x"00",x"00",x"00",x"7E",x"02",x"02",x"02",x"1A",x"26",x"40",x"40",x"42",x"22",x"1C",x"00",x"00"), --! "5",21*/
  (x"00",x"00",x"00",x"38",x"24",x"02",x"02",x"1A",x"26",x"42",x"42",x"42",x"24",x"18",x"00",x"00"), --! "6",22*/
  (x"00",x"00",x"00",x"7E",x"22",x"22",x"10",x"10",x"08",x"08",x"08",x"08",x"08",x"08",x"00",x"00"), --! "7",23*/
  (x"00",x"00",x"00",x"3C",x"42",x"42",x"42",x"24",x"18",x"24",x"42",x"42",x"42",x"3C",x"00",x"00"), --! "8",24*/
  (x"00",x"00",x"00",x"18",x"24",x"42",x"42",x"42",x"64",x"58",x"40",x"40",x"24",x"1C",x"00",x"00"), --! "9",25*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00"), --! ":",26*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"04"), --! ";",27*/
  (x"00",x"00",x"00",x"40",x"20",x"10",x"08",x"04",x"02",x"04",x"08",x"10",x"20",x"40",x"00",x"00"), --! "<",28*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"7F",x"00",x"00",x"00",x"7F",x"00",x"00",x"00",x"00",x"00"), --! "=",29*/
  (x"00",x"00",x"00",x"02",x"04",x"08",x"10",x"20",x"40",x"20",x"10",x"08",x"04",x"02",x"00",x"00"), --! ">",30*/
  (x"00",x"00",x"00",x"3C",x"42",x"42",x"46",x"40",x"20",x"10",x"10",x"00",x"18",x"18",x"00",x"00"), --! "?",31*/
  (x"00",x"00",x"00",x"1C",x"22",x"5A",x"55",x"55",x"55",x"55",x"2D",x"42",x"22",x"1C",x"00",x"00"), --! "@",32*/
  (x"00",x"00",x"00",x"08",x"08",x"18",x"14",x"14",x"24",x"3C",x"22",x"42",x"42",x"E7",x"00",x"00"), --! "A",33*/
  (x"00",x"00",x"00",x"1F",x"22",x"22",x"22",x"1E",x"22",x"42",x"42",x"42",x"22",x"1F",x"00",x"00"), --! "B",34*/
  (x"00",x"00",x"00",x"7C",x"42",x"42",x"01",x"01",x"01",x"01",x"01",x"42",x"22",x"1C",x"00",x"00"), --! "C",35*/
  (x"00",x"00",x"00",x"1F",x"22",x"42",x"42",x"42",x"42",x"42",x"42",x"42",x"22",x"1F",x"00",x"00"), --! "D",36*/
  (x"00",x"00",x"00",x"3F",x"42",x"12",x"12",x"1E",x"12",x"12",x"02",x"42",x"42",x"3F",x"00",x"00"), --! "E",37*/
  (x"00",x"00",x"00",x"3F",x"42",x"12",x"12",x"1E",x"12",x"12",x"02",x"02",x"02",x"07",x"00",x"00"), --! "F",38*/
  (x"00",x"00",x"00",x"3C",x"22",x"22",x"01",x"01",x"01",x"71",x"21",x"22",x"22",x"1C",x"00",x"00"), --! "G",39*/
  (x"00",x"00",x"00",x"E7",x"42",x"42",x"42",x"42",x"7E",x"42",x"42",x"42",x"42",x"E7",x"00",x"00"), --! "H",40*/
  (x"00",x"00",x"00",x"3E",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"3E",x"00",x"00"), --! "I",41*/
  (x"00",x"00",x"00",x"7C",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"11",x"0F"), --! "J",42*/
  (x"00",x"00",x"00",x"77",x"22",x"12",x"0A",x"0E",x"0A",x"12",x"12",x"22",x"22",x"77",x"00",x"00"), --! "K",43*/
  (x"00",x"00",x"00",x"07",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"42",x"7F",x"00",x"00"), --! "L",44*/
  (x"00",x"00",x"00",x"77",x"36",x"36",x"36",x"36",x"2A",x"2A",x"2A",x"2A",x"2A",x"6B",x"00",x"00"), --! "M",45*/
  (x"00",x"00",x"00",x"E3",x"46",x"46",x"4A",x"4A",x"52",x"52",x"52",x"62",x"62",x"47",x"00",x"00"), --! "N",46*/
  (x"00",x"00",x"00",x"1C",x"22",x"41",x"41",x"41",x"41",x"41",x"41",x"41",x"22",x"1C",x"00",x"00"), --! "O",47*/
  (x"00",x"00",x"00",x"3F",x"42",x"42",x"42",x"42",x"3E",x"02",x"02",x"02",x"02",x"07",x"00",x"00"), --! "P",48*/
  (x"00",x"00",x"00",x"1C",x"22",x"41",x"41",x"41",x"41",x"41",x"4D",x"53",x"32",x"1C",x"60",x"00"), --! "Q",49*/
  (x"00",x"00",x"00",x"3F",x"42",x"42",x"42",x"3E",x"12",x"12",x"22",x"22",x"42",x"C7",x"00",x"00"), --! "R",50*/
  (x"00",x"00",x"00",x"7C",x"42",x"42",x"02",x"04",x"18",x"20",x"40",x"42",x"42",x"3E",x"00",x"00"), --! "S",51*/
  (x"00",x"00",x"00",x"7F",x"49",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"1C",x"00",x"00"), --! "T",52*/
  (x"00",x"00",x"00",x"E7",x"42",x"42",x"42",x"42",x"42",x"42",x"42",x"42",x"42",x"3C",x"00",x"00"), --! "U",53*/
  (x"00",x"00",x"00",x"E7",x"42",x"42",x"22",x"24",x"24",x"14",x"14",x"18",x"08",x"08",x"00",x"00"), --! "V",54*/
  (x"00",x"00",x"00",x"6B",x"49",x"49",x"49",x"49",x"55",x"55",x"36",x"22",x"22",x"22",x"00",x"00"), --! "W",55*/
  (x"00",x"00",x"00",x"E7",x"42",x"24",x"24",x"18",x"18",x"18",x"24",x"24",x"42",x"E7",x"00",x"00"), --! "X",56*/
  (x"00",x"00",x"00",x"77",x"22",x"22",x"14",x"14",x"08",x"08",x"08",x"08",x"08",x"1C",x"00",x"00"), --! "Y",57*/
  (x"00",x"00",x"00",x"7E",x"21",x"20",x"10",x"10",x"08",x"04",x"04",x"42",x"42",x"3F",x"00",x"00"), --! "Z",58*/
  (x"00",x"78",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"78",x"00"), --! "[",59*/
  (x"00",x"00",x"02",x"02",x"04",x"04",x"08",x"08",x"08",x"10",x"10",x"20",x"20",x"20",x"40",x"40"), --! "\",60*/
  (x"00",x"1E",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"1E",x"00"), --! "]",61*/
  (x"00",x"38",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"), --! "^",62*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF"), --! "_",63*/
  (x"00",x"06",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"), --! "`",64*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"42",x"78",x"44",x"42",x"42",x"FC",x"00",x"00"), --! "a",65*/
  (x"00",x"00",x"00",x"03",x"02",x"02",x"02",x"1A",x"26",x"42",x"42",x"42",x"26",x"1A",x"00",x"00"), --! "b",66*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"44",x"02",x"02",x"02",x"44",x"38",x"00",x"00"), --! "c",67*/
  (x"00",x"00",x"00",x"60",x"40",x"40",x"40",x"78",x"44",x"42",x"42",x"42",x"64",x"D8",x"00",x"00"), --! "d",68*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"42",x"7E",x"02",x"02",x"42",x"3C",x"00",x"00"), --! "e",69*/
  (x"00",x"00",x"00",x"F0",x"88",x"08",x"08",x"7E",x"08",x"08",x"08",x"08",x"08",x"3E",x"00",x"00"), --! "f",70*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"22",x"22",x"1C",x"02",x"3C",x"42",x"42",x"3C"), --! "g",71*/
  (x"00",x"00",x"00",x"03",x"02",x"02",x"02",x"3A",x"46",x"42",x"42",x"42",x"42",x"E7",x"00",x"00"), --! "h",72*/
  (x"00",x"00",x"00",x"0C",x"0C",x"00",x"00",x"0E",x"08",x"08",x"08",x"08",x"08",x"3E",x"00",x"00"), --! "i",73*/
  (x"00",x"00",x"00",x"30",x"30",x"00",x"00",x"38",x"20",x"20",x"20",x"20",x"20",x"20",x"22",x"1E"), --! "j",74*/
  (x"00",x"00",x"00",x"03",x"02",x"02",x"02",x"72",x"12",x"0A",x"16",x"12",x"22",x"77",x"00",x"00"), --! "k",75*/
  (x"00",x"00",x"00",x"0E",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"3E",x"00",x"00"), --! "l",76*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7F",x"92",x"92",x"92",x"92",x"92",x"B7",x"00",x"00"), --! "m",77*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3B",x"46",x"42",x"42",x"42",x"42",x"E7",x"00",x"00"), --! "n",78*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3C",x"42",x"42",x"42",x"42",x"42",x"3C",x"00",x"00"), --! "o",79*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"1B",x"26",x"42",x"42",x"42",x"22",x"1E",x"02",x"07"), --! "p",80*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"78",x"44",x"42",x"42",x"42",x"44",x"78",x"40",x"E0"), --! "q",81*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"77",x"4C",x"04",x"04",x"04",x"04",x"1F",x"00",x"00"), --! "r",82*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"42",x"02",x"3C",x"40",x"42",x"3E",x"00",x"00"), --! "s",83*/
  (x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"3E",x"08",x"08",x"08",x"08",x"08",x"30",x"00",x"00"), --! "t",84*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"63",x"42",x"42",x"42",x"42",x"62",x"DC",x"00",x"00"), --! "u",85*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E7",x"42",x"24",x"24",x"14",x"08",x"08",x"00",x"00"), --! "v",86*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EB",x"49",x"49",x"55",x"55",x"22",x"22",x"00",x"00"), --! "w",87*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"76",x"24",x"18",x"18",x"18",x"24",x"6E",x"00",x"00"), --! "x",88*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E7",x"42",x"24",x"24",x"14",x"18",x"08",x"08",x"07"), --! "y",89*/
  (x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7E",x"22",x"10",x"08",x"08",x"44",x"7E",x"00",x"00"), --! "z",90*/
  (x"00",x"C0",x"20",x"20",x"20",x"20",x"20",x"10",x"20",x"20",x"20",x"20",x"20",x"20",x"C0",x"00"), --! "{",91*/
  (x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10"), --! "|",92*/
  (x"00",x"06",x"08",x"08",x"08",x"08",x"08",x"10",x"08",x"08",x"08",x"08",x"08",x"08",x"06",x"00"), --! "}",93*/
  (x"0C",x"32",x"C2",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")  --! "~",94*/
  );


end package ascii_pkg;
-------------------------------------------------------------------------------
package body ascii_pkg is

end package body ascii_pkg;