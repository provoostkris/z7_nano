library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-------------------------------------------------------------------------------
package pmod_lcd_pkg is

  -- factor for the clock divider , to reduce the SPI clock from the system clock
  constant c_clk_reduce             : integer := 2;
  -- proper reset time
  -- 1 clk = 20 ns ==> 1 us = 50x
  -- and divide by the clock reduction factor
  constant c_rst_time_act           : integer :=    1000 * 50 / 2**(c_clk_reduce+1); -- minimum   1_000 us
  constant c_rst_time_hld           : integer := 200_000 * 50 / 2**(c_clk_reduce+1); -- minimum 200_000 us
  constant c_sleep_out              : integer := 150_000 * 50 / 2**(c_clk_reduce+1); -- minimum 150_000 us

  -- constants found in the LCD controller datasheet
  constant c_bits_565         : integer := 5+6+5;
  constant c_bits_666         : integer := 8+8+8;
  constant c_bits             : integer := c_bits_565;
  constant c_hori             : integer := 160;   --! Horizontal amount of pixels
  constant c_vert             : integer := 80;    --! Vertical amount of pixels
  constant c_pixl             : integer := c_hori * c_vert;  --! total amount of pixels

  constant c_off_h            : integer := 2;   --! offset to 1st pixel in hori
  constant c_off_v            : integer := 27;  --! offset to 1st pixel in vert

  constant c_SLPOUT           : std_logic_vector(7 downto 0) := x"11";  --! sleep out
  constant c_DISPOFF          : std_logic_vector(7 downto 0) := x"28";  --! display off
  constant c_DISPON           : std_logic_vector(7 downto 0) := x"29";  --! display on
  constant c_CASET            : std_logic_vector(7 downto 0) := x"2A";  --! column address set
  constant c_RASET            : std_logic_vector(7 downto 0) := x"2B";  --! row address set
  constant c_RAMWR            : std_logic_vector(7 downto 0) := x"2C";  --! RAM write
  constant c_MADCTL           : std_logic_vector(7 downto 0) := x"36";  --! axis control
  constant c_COLMOD           : std_logic_vector(7 downto 0) := x"3A";  --! color mode

  -- just some random values to driver the display for testing
  constant c_tst_colors       : std_logic_vector(24-1 downto 0) :=  "00001111" &
                                                                    "11001100" &
                                                                    "00110011" ;

  -- create arrays for pixel map stores
  type t_raw_arr  is array (integer range <>) of std_logic_vector(24-1 downto 0); -- raw pixel map
  type t_rgb_arr  is array (integer range <>) of integer range 0 to 255;              -- rgb array
  type t_clr_arr  is array (integer range <>) of t_rgb_arr( 0 to 2);                  -- color array
  type t_cnt_arr  is array (integer range <>) of integer range 0 to c_bits-1;         -- counter array

  constant c_color_map : t_clr_arr( 0 to c_pixl-1) :=
  -- manually modified the first three pixels to be fixed for r & g & b to check the timing and alignment
((255, 127, 127), (127, 127, 127), (255, 0, 255), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 1, 3), (0, 0, 2), (0, 0, 0), (2, 0, 0), (2, 0, 0), (2, 0, 0), (0, 0, 2), (0, 0, 6), (205, 212, 223), (203, 212, 227), (202, 213, 231), (201, 213, 233), (203, 214, 234), (205, 215, 234), (206, 214, 233), (207, 214, 232), (210, 216, 234), (207, 216, 233), (201, 219, 233), (201, 220, 234), (203, 219, 234), (206, 216, 233), (213, 216, 235), (216, 217, 237), (208, 215, 234), (210, 221, 239), (208, 224, 240), (208, 224, 240), (209, 222, 239), (210, 221, 239), (213, 224, 242), (212, 220, 241), (220, 221, 247), (219, 221, 243), (216, 226, 234), (222, 233, 238), (219, 226, 237), (221, 227, 243), (214, 227, 243), (214, 229, 241), (214, 229, 231), (220, 239, 236), (210, 236, 234), (210, 235, 238), (217, 230, 244), (227, 234, 251), (223, 230, 241), (226, 233, 243), (226, 235, 248), (224, 229, 244), (228, 224, 240), (232, 227, 239), (238, 239, 242), (224, 234, 236), (215, 235, 245), (216, 238, 254), (223, 237, 255), (221, 229, 249), (232, 237, 249), (233, 235, 244), (228, 228, 242), (235, 237, 250), (227, 236, 243), (228, 239, 244), (228, 237, 243), (233, 242, 247), (234, 244, 245), (229, 239, 240), (230, 239, 247), (230, 238, 251), (228, 235, 251), (233, 240, 255), (233, 240, 249), (234, 240, 247), (235, 241, 248), (236, 240, 251), (238, 240, 255), (239, 239, 255), (239, 239, 253), (238, 239, 250), (239, 240, 250), (239, 242, 251), (239, 241, 252), (239, 241, 253), (239, 241, 253), (240, 241, 252), (240, 241, 250), (241, 242, 248), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 1, 2), (0, 1, 2), (0, 0, 0), (2, 0, 0), (2, 0, 0), (2, 0, 0), (0, 0, 2), (0, 0, 6), (205, 212, 223), (203, 212, 227), (201, 214, 231), (201, 214, 233), (202, 214, 234), (205, 215, 234), (206, 215, 232), (207, 214, 231), (208, 215, 232), (205, 215, 231), (203, 218, 233), (203, 219, 234), (204, 219, 234), (205, 216, 233), (210, 216, 234), (212, 217, 236), (212, 220, 239), (207, 217, 235), (203, 216, 232), (208, 221, 237), (212, 222, 238), (216, 224, 239), (216, 222, 238), (221, 225, 243), (217, 221, 242), (216, 220, 239), (216, 224, 235), (215, 225, 233), (216, 227, 239), (215, 227, 242), (218, 231, 247), (220, 232, 245), (219, 230, 235), (217, 230, 231), (210, 230, 231), (217, 236, 242), (218, 231, 245), (225, 234, 249), (224, 231, 242), (224, 231, 241), (223, 231, 242), (231, 231, 242), (245, 226, 239), (253, 222, 234), (239, 203, 211), (250, 221, 230), (239, 230, 244), (228, 231, 250), (224, 231, 253), (233, 241, 255), (230, 234, 245), (227, 230, 238), (235, 239, 249), (225, 230, 240), (228, 236, 242), (227, 236, 241), (225, 234, 241), (225, 234, 240), (226, 236, 237), (227, 237, 238), (232, 241, 248), (234, 242, 253), (230, 238, 252), (231, 239, 252), (233, 240, 249), (234, 240, 247), (235, 241, 248), (236, 240, 250), (237, 239, 253), (239, 240, 254), (238, 239, 251), (238, 239, 249), (239, 241, 250), (238, 241, 250), (239, 241, 252), (239, 241, 253), (239, 241, 253), (240, 241, 252), (240, 241, 250), (241, 242, 248), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 1, 2), (0, 1, 1), (0, 0, 0), (2, 0, 0), (2, 0, 0), (2, 0, 0), (0, 0, 2), (0, 0, 6), (205, 212, 223), (202, 213, 227), (201, 214, 231), (200, 214, 233), (202, 215, 233), (204, 215, 233), (205, 215, 231), (205, 215, 230), (204, 216, 230), (204, 216, 231), (206, 216, 232), (208, 218, 235), (206, 219, 236), (205, 218, 235), (204, 218, 235), (206, 219, 236), (211, 221, 239), (210, 218, 236), (214, 221, 237), (220, 226, 240), (215, 220, 232), (218, 221, 231), (206, 203, 213), (205, 205, 215), (214, 222, 234), (215, 226, 238), (220, 225, 240), (218, 226, 241), (212, 231, 245), (210, 231, 245), (215, 228, 243), (221, 228, 243), (225, 227, 240), (224, 226, 237), (224, 229, 240), (226, 236, 246), (215, 229, 240), (218, 230, 243), (224, 230, 244), (226, 230, 241), (223, 231, 235), (233, 224, 227), (255, 210, 216), (232, 150, 161), (206, 96, 113), (211, 106, 127), (255, 189, 213), (255, 228, 252), (231, 224, 247), (215, 221, 239), (226, 230, 240), (229, 234, 239), (226, 236, 239), (232, 243, 246), (228, 236, 240), (231, 239, 244), (234, 242, 251), (231, 240, 247), (230, 240, 242), (231, 241, 242), (230, 239, 243), (229, 238, 244), (231, 239, 249), (233, 241, 251), (233, 240, 248), (234, 240, 247), (235, 241, 247), (236, 241, 247), (237, 240, 248), (238, 240, 248), (238, 240, 247), (238, 239, 247), (238, 240, 248), (237, 240, 249), (238, 240, 251), (238, 240, 252), (239, 241, 253), (240, 241, 252), (240, 241, 250), (241, 242, 248), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 1), (0, 1, 1), (0, 0, 0), (2, 0, 0), (2, 0, 0), (2, 0, 0), (0, 0, 2), (0, 1, 6), (204, 212, 223), (201, 213, 227), (200, 214, 231), (199, 214, 232), (201, 215, 233), (203, 216, 233), (205, 215, 231), (204, 216, 230), (202, 219, 231), (202, 218, 231), (208, 217, 233), (210, 217, 234), (207, 218, 235), (205, 220, 235), (202, 221, 235), (203, 222, 236), (205, 219, 235), (213, 222, 238), (217, 222, 236), (211, 213, 225), (200, 202, 210), (219, 217, 223), (212, 204, 210), (214, 209, 214), (215, 223, 227), (218, 229, 237), (219, 222, 237), (221, 228, 245), (207, 229, 242), (212, 234, 246), (214, 225, 237), (224, 226, 238), (220, 217, 228), (228, 223, 235), (229, 228, 241), (226, 230, 242), (218, 229, 240), (221, 233, 244), (226, 233, 244), (225, 229, 238), (223, 230, 232), (251, 231, 233), (237, 163, 169), (209, 90, 103), (230, 74, 97), (210, 55, 86), (171, 57, 92), (229, 156, 192), (253, 221, 253), (215, 205, 232), (238, 231, 249), (229, 227, 239), (228, 232, 239), (226, 234, 239), (226, 235, 243), (226, 234, 245), (225, 233, 246), (226, 234, 246), (228, 237, 243), (233, 243, 245), (233, 243, 244), (229, 238, 242), (230, 239, 246), (231, 238, 247), (233, 240, 249), (234, 240, 248), (235, 241, 247), (236, 241, 245), (237, 241, 245), (237, 240, 245), (238, 240, 245), (238, 240, 247), (237, 240, 248), (237, 240, 249), (237, 239, 250), (238, 240, 252), (238, 240, 252), (240, 241, 252), (240, 241, 250), (241, 242, 248), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (1, 0, 0), (2, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 2), (0, 1, 6), (203, 213, 223), (200, 213, 227), (199, 215, 230), (199, 215, 232), (200, 216, 233), (203, 216, 233), (205, 216, 231), (203, 217, 230), (199, 222, 232), (199, 221, 232), (206, 218, 231), (207, 216, 230), (206, 217, 230), (203, 219, 231), (201, 224, 233), (201, 225, 235), (204, 222, 233), (210, 222, 234), (212, 219, 230), (208, 209, 218), (200, 199, 205), (224, 219, 223), (223, 212, 215), (230, 221, 223), (222, 222, 224), (219, 224, 228), (217, 221, 232), (216, 225, 238), (211, 228, 238), (214, 231, 239), (222, 228, 234), (230, 229, 233), (228, 220, 224), (233, 226, 232), (227, 227, 235), (221, 225, 235), (226, 233, 243), (224, 232, 241), (220, 229, 235), (221, 228, 232), (221, 223, 229), (255, 224, 231), (248, 152, 163), (231, 88, 106), (216, 40, 69), (193, 17, 56), (188, 42, 90), (197, 87, 139), (255, 195, 246), (255, 220, 255), (254, 224, 255), (254, 234, 255), (247, 233, 254), (236, 232, 249), (235, 245, 255), (234, 248, 255), (228, 237, 255), (230, 237, 255), (223, 231, 241), (227, 236, 240), (232, 242, 242), (231, 241, 241), (234, 242, 247), (230, 237, 246), (233, 240, 251), (234, 239, 250), (234, 240, 247), (236, 241, 246), (237, 241, 244), (237, 241, 244), (237, 240, 246), (237, 240, 247), (236, 239, 247), (237, 240, 249), (237, 239, 250), (237, 239, 251), (238, 240, 252), (240, 241, 252), (240, 241, 250), (242, 243, 249), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (1, 0, 0), (2, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 3), (0, 1, 7), (203, 213, 223), (200, 214, 227), (199, 215, 230), (198, 215, 231), (200, 216, 232), (202, 216, 232), (205, 216, 230), (203, 217, 230), (197, 221, 231), (197, 221, 231), (204, 218, 230), (205, 215, 227), (205, 215, 226), (205, 218, 228), (203, 223, 231), (203, 225, 232), (205, 225, 233), (207, 222, 230), (214, 221, 230), (223, 223, 231), (224, 217, 223), (234, 223, 227), (227, 212, 215), (230, 217, 219), (229, 221, 224), (219, 215, 220), (225, 222, 231), (223, 224, 234), (224, 231, 239), (218, 226, 230), (225, 228, 227), (226, 224, 220), (234, 225, 220), (236, 228, 226), (229, 230, 234), (221, 226, 234), (225, 230, 241), (224, 228, 236), (230, 231, 232), (244, 233, 232), (255, 226, 230), (255, 192, 201), (255, 128, 141), (242, 67, 89), (213, 22, 56), (189, 0, 47), (223, 56, 118), (219, 81, 151), (185, 82, 156), (185, 109, 181), (189, 130, 195), (219, 171, 228), (233, 191, 238), (229, 201, 242), (193, 186, 227), (143, 147, 185), (223, 228, 255), (237, 243, 255), (230, 238, 250), (227, 236, 240), (230, 240, 239), (231, 240, 240), (235, 242, 249), (233, 240, 251), (234, 239, 253), (234, 239, 252), (235, 239, 249), (236, 241, 247), (237, 241, 245), (237, 240, 245), (237, 240, 247), (237, 240, 249), (237, 240, 249), (237, 240, 249), (237, 239, 250), (237, 239, 251), (238, 240, 252), (240, 241, 252), (240, 241, 250), (242, 243, 249), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (1, 0, 0), (1, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 3), (0, 1, 7), (203, 213, 223), (200, 214, 227), (199, 215, 230), (198, 215, 231), (200, 216, 231), (202, 217, 231), (205, 216, 229), (203, 216, 230), (198, 217, 231), (199, 220, 232), (202, 219, 230), (203, 215, 226), (207, 214, 224), (210, 217, 226), (209, 219, 226), (207, 222, 227), (206, 225, 230), (206, 222, 228), (211, 218, 225), (224, 221, 229), (230, 217, 225), (236, 216, 223), (236, 215, 220), (239, 220, 225), (234, 220, 228), (223, 209, 218), (226, 209, 217), (238, 223, 229), (226, 217, 221), (224, 220, 220), (220, 221, 213), (220, 219, 206), (221, 210, 196), (224, 214, 204), (227, 227, 226), (220, 226, 232), (220, 228, 238), (231, 231, 238), (246, 228, 225), (252, 201, 196), (248, 149, 150), (204, 57, 64), (218, 22, 35), (237, 22, 46), (238, 35, 72), (238, 48, 102), (190, 14, 89), (204, 47, 137), (141, 6, 108), (129, 15, 121), (138, 43, 147), (134, 50, 147), (118, 37, 123), (105, 38, 117), (113, 71, 148), (92, 70, 136), (187, 182, 228), (223, 228, 255), (233, 241, 254), (233, 242, 246), (235, 244, 244), (230, 238, 241), (232, 239, 249), (231, 236, 251), (233, 238, 253), (235, 238, 253), (235, 239, 251), (236, 240, 251), (237, 240, 250), (237, 239, 250), (237, 239, 251), (237, 239, 251), (237, 240, 249), (237, 240, 249), (237, 239, 250), (237, 239, 251), (238, 240, 252), (240, 241, 252), (240, 241, 250), (242, 243, 249), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 4), (0, 1, 8), (203, 213, 223), (200, 214, 227), (199, 215, 230), (198, 215, 231), (200, 216, 231), (203, 217, 231), (205, 216, 229), (204, 216, 229), (201, 215, 231), (202, 218, 234), (203, 218, 231), (204, 216, 228), (209, 214, 226), (214, 217, 227), (214, 218, 228), (210, 218, 227), (206, 221, 227), (211, 226, 232), (215, 221, 228), (219, 214, 221), (226, 206, 213), (233, 203, 209), (242, 209, 212), (242, 210, 214), (242, 215, 224), (228, 201, 210), (219, 184, 190), (247, 211, 214), (217, 188, 190), (233, 212, 210), (223, 212, 201), (229, 220, 204), (216, 203, 184), (217, 205, 191), (229, 225, 223), (224, 225, 231), (222, 228, 236), (240, 231, 234), (243, 200, 193), (212, 122, 112), (209, 63, 57), (214, 23, 24), (235, 11, 21), (228, 0, 22), (214, 13, 50), (203, 20, 75), (185, 11, 88), (174, 11, 107), (157, 6, 118), (170, 35, 156), (113, 0, 119), (142, 36, 156), (78, 0, 90), (100, 13, 117), (150, 79, 184), (199, 152, 240), (187, 174, 228), (223, 228, 255), (230, 238, 249), (225, 235, 237), (231, 239, 240), (230, 238, 242), (234, 239, 252), (233, 238, 253), (234, 237, 252), (235, 239, 252), (235, 239, 251), (236, 239, 252), (237, 239, 253), (237, 239, 253), (237, 239, 252), (237, 239, 251), (238, 241, 250), (237, 240, 249), (237, 239, 250), (238, 240, 252), (238, 240, 252), (240, 241, 252), (240, 241, 250), (242, 243, 249), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 4), (0, 1, 8), (205, 215, 225), (200, 214, 227), (197, 213, 228), (199, 215, 231), (201, 216, 231), (202, 215, 229), (205, 216, 228), (207, 216, 230), (206, 214, 233), (207, 217, 236), (205, 218, 234), (206, 217, 231), (207, 212, 227), (212, 213, 228), (216, 216, 232), (214, 217, 232), (209, 218, 231), (211, 221, 231), (216, 219, 227), (234, 225, 230), (216, 190, 193), (195, 154, 154), (219, 168, 165), (230, 178, 176), (241, 197, 202), (246, 201, 207), (200, 141, 145), (242, 182, 184), (242, 191, 190), (243, 201, 197), (230, 197, 188), (237, 214, 199), (220, 205, 186), (224, 212, 199), (242, 227, 230), (235, 225, 233), (227, 228, 231), (247, 226, 222), (242, 167, 155), (219, 93, 78), (232, 58, 46), (227, 21, 15), (229, 8, 11), (215, 0, 16), (191, 5, 37), (179, 11, 61), (204, 43, 111), (187, 32, 117), (161, 11, 115), (163, 21, 139), (175, 46, 173), (178, 65, 192), (99, 3, 121), (98, 8, 125), (112, 17, 142), (158, 85, 190), (191, 170, 227), (203, 209, 233), (231, 240, 247), (223, 233, 232), (233, 241, 242), (235, 241, 246), (232, 237, 250), (233, 236, 251), (232, 236, 247), (238, 242, 251), (235, 238, 248), (235, 237, 249), (236, 238, 254), (235, 237, 252), (237, 239, 250), (238, 241, 250), (237, 240, 249), (237, 240, 249), (237, 239, 250), (238, 240, 252), (238, 240, 252), (239, 240, 251), (240, 241, 250), (241, 242, 248), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 4), (0, 1, 8), (202, 212, 222), (199, 212, 225), (198, 214, 229), (200, 216, 232), (204, 218, 234), (208, 220, 234), (206, 217, 228), (204, 212, 225), (208, 215, 233), (211, 219, 239), (205, 215, 232), (213, 223, 239), (210, 216, 233), (213, 217, 235), (207, 210, 229), (215, 219, 238), (214, 223, 240), (212, 221, 235), (214, 218, 226), (230, 222, 225), (221, 194, 192), (201, 156, 149), (237, 175, 164), (251, 183, 173), (246, 181, 175), (225, 154, 151), (233, 148, 145), (255, 171, 168), (255, 190, 185), (194, 124, 117), (207, 147, 137), (236, 191, 178), (240, 211, 195), (233, 212, 201), (212, 186, 189), (221, 199, 203), (234, 225, 218), (229, 194, 178), (242, 143, 121), (255, 106, 85), (242, 50, 36), (228, 16, 10), (225, 12, 16), (206, 9, 26), (158, 0, 27), (142, 0, 46), (150, 16, 76), (142, 13, 87), (126, 0, 87), (138, 7, 116), (145, 18, 142), (176, 61, 189), (118, 27, 146), (82, 0, 115), (103, 2, 131), (136, 56, 163), (177, 154, 207), (216, 223, 242), (226, 235, 241), (236, 246, 246), (233, 241, 244), (229, 235, 242), (225, 230, 243), (240, 244, 255), (241, 245, 253), (231, 236, 241), (236, 239, 246), (238, 240, 251), (235, 237, 252), (233, 235, 249), (240, 243, 251), (235, 238, 244), (237, 240, 248), (237, 240, 249), (237, 239, 250), (237, 239, 251), (238, 240, 252), (239, 240, 251), (239, 240, 249), (240, 241, 247), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 4), (0, 1, 8), (203, 213, 223), (203, 216, 229), (202, 217, 232), (199, 214, 230), (198, 211, 226), (202, 213, 226), (203, 211, 222), (201, 209, 221), (202, 211, 227), (206, 216, 233), (209, 218, 235), (201, 211, 228), (203, 214, 231), (213, 226, 244), (204, 217, 237), (209, 223, 243), (207, 221, 241), (211, 224, 239), (216, 226, 233), (226, 225, 224), (232, 212, 202), (240, 199, 182), (238, 171, 152), (217, 134, 112), (242, 152, 129), (207, 106, 85), (226, 111, 96), (244, 125, 112), (230, 118, 105), (160, 57, 44), (206, 114, 101), (255, 181, 168), (255, 216, 204), (255, 218, 210), (213, 173, 172), (233, 200, 194), (255, 237, 213), (238, 188, 154), (247, 133, 97), (255, 99, 69), (254, 56, 45), (223, 12, 14), (209, 7, 21), (193, 18, 42), (134, 2, 36), (102, 0, 41), (76, 0, 38), (71, 0, 47), (81, 0, 66), (110, 6, 102), (142, 26, 141), (182, 73, 193), (92, 8, 120), (59, 0, 93), (88, 0, 115), (123, 54, 147), (190, 172, 215), (239, 247, 255), (221, 230, 236), (218, 227, 232), (227, 234, 242), (243, 249, 255), (236, 241, 254), (234, 238, 248), (232, 236, 240), (238, 242, 244), (234, 237, 242), (240, 243, 251), (235, 237, 249), (240, 243, 253), (233, 237, 240), (243, 247, 250), (237, 240, 247), (237, 240, 249), (237, 239, 250), (237, 239, 251), (237, 239, 251), (239, 240, 251), (239, 240, 249), (240, 241, 247), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 4), (0, 1, 8), (203, 213, 223), (202, 214, 227), (200, 214, 230), (200, 213, 230), (201, 213, 228), (205, 214, 228), (208, 215, 226), (209, 216, 227), (209, 217, 229), (212, 220, 233), (202, 205, 220), (215, 218, 233), (213, 219, 234), (203, 213, 229), (209, 223, 241), (204, 220, 238), (207, 223, 241), (208, 224, 238), (214, 228, 235), (221, 226, 223), (234, 222, 209), (255, 228, 209), (218, 156, 134), (170, 85, 57), (228, 123, 87), (214, 90, 55), (225, 82, 57), (253, 105, 85), (232, 94, 75), (194, 66, 48), (207, 88, 73), (218, 113, 102), (205, 116, 110), (243, 168, 164), (235, 171, 168), (229, 177, 164), (235, 193, 162), (245, 179, 138), (255, 135, 96), (249, 74, 45), (250, 45, 35), (220, 9, 15), (194, 3, 20), (164, 8, 35), (106, 0, 35), (67, 0, 33), (68, 0, 51), (92, 11, 86), (103, 11, 101), (107, 2, 107), (145, 26, 146), (140, 26, 149), (100, 7, 122), (81, 0, 107), (99, 7, 117), (155, 85, 171), (241, 223, 255), (224, 232, 245), (230, 238, 252), (226, 233, 249), (235, 241, 255), (212, 216, 234), (213, 216, 231), (237, 241, 252), (239, 242, 248), (242, 246, 249), (232, 235, 241), (174, 177, 185), (232, 235, 243), (233, 236, 243), (243, 247, 249), (232, 236, 238), (236, 239, 246), (237, 240, 249), (237, 239, 250), (237, 239, 251), (237, 239, 251), (238, 239, 250), (238, 239, 248), (239, 240, 246), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 4), (0, 1, 8), (204, 212, 223), (200, 211, 225), (198, 211, 227), (200, 213, 230), (205, 215, 231), (207, 215, 229), (208, 213, 225), (208, 212, 222), (207, 212, 219), (201, 203, 210), (210, 204, 213), (222, 213, 223), (212, 206, 215), (223, 222, 231), (212, 218, 230), (206, 217, 230), (208, 223, 237), (206, 222, 234), (211, 227, 233), (217, 226, 225), (226, 220, 211), (245, 220, 206), (245, 198, 180), (241, 164, 137), (247, 137, 92), (187, 46, 0), (208, 39, 6), (232, 57, 31), (227, 69, 43), (212, 66, 43), (249, 109, 92), (203, 65, 56), (173, 36, 36), (207, 83, 85), (228, 129, 124), (226, 147, 131), (230, 165, 134), (255, 169, 133), (255, 116, 86), (238, 51, 31), (227, 13, 5), (217, 5, 9), (185, 4, 19), (135, 0, 20), (89, 4, 36), (59, 0, 41), (108, 15, 98), (153, 41, 149), (165, 39, 164), (160, 27, 163), (163, 26, 166), (121, 0, 127), (108, 0, 120), (166, 57, 176), (148, 37, 148), (163, 81, 164), (238, 216, 252), (227, 234, 252), (232, 237, 255), (230, 234, 255), (222, 225, 255), (122, 124, 154), (194, 196, 216), (235, 237, 251), (235, 237, 249), (226, 228, 240), (213, 215, 227), (228, 231, 240), (239, 242, 249), (243, 246, 251), (230, 234, 237), (237, 240, 245), (236, 239, 247), (236, 239, 248), (237, 239, 250), (237, 239, 251), (237, 239, 251), (238, 239, 250), (238, 239, 248), (239, 240, 246), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 4), (0, 1, 8), (204, 212, 223), (203, 214, 227), (202, 214, 230), (201, 212, 229), (201, 210, 225), (204, 210, 224), (209, 213, 225), (215, 215, 224), (216, 213, 217), (197, 188, 191), (224, 205, 209), (218, 194, 198), (226, 201, 205), (226, 205, 209), (227, 215, 220), (221, 218, 226), (219, 225, 234), (211, 222, 231), (205, 217, 224), (217, 225, 229), (233, 229, 228), (222, 204, 200), (246, 212, 204), (241, 177, 156), (217, 109, 63), (255, 108, 57), (250, 68, 31), (223, 35, 6), (192, 27, 0), (249, 93, 71), (255, 119, 109), (255, 101, 101), (240, 63, 71), (220, 55, 62), (209, 73, 73), (215, 102, 93), (237, 141, 123), (254, 141, 123), (238, 74, 64), (215, 17, 14), (215, 0, 3), (224, 12, 25), (198, 11, 36), (136, 0, 23), (85, 0, 31), (62, 0, 42), (115, 9, 102), (144, 20, 141), (142, 12, 148), (168, 33, 178), (184, 46, 190), (150, 12, 153), (181, 46, 182), (191, 64, 189), (188, 70, 181), (243, 160, 241), (253, 230, 255), (233, 239, 255), (196, 199, 244), (181, 182, 237), (155, 155, 207), (174, 174, 216), (210, 210, 236), (231, 232, 251), (226, 227, 248), (215, 216, 237), (219, 220, 239), (243, 245, 255), (211, 214, 220), (227, 231, 235), (242, 245, 252), (234, 237, 246), (237, 240, 249), (237, 240, 249), (237, 239, 250), (237, 239, 251), (237, 239, 251), (238, 239, 250), (238, 239, 248), (239, 240, 246), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 4), (0, 1, 8), (201, 209, 220), (204, 214, 229), (204, 215, 232), (202, 212, 229), (204, 211, 227), (211, 216, 229), (212, 214, 226), (212, 208, 216), (230, 214, 217), (223, 197, 197), (221, 185, 185), (235, 191, 190), (254, 203, 201), (211, 161, 160), (238, 198, 197), (234, 208, 209), (220, 211, 214), (225, 225, 232), (221, 224, 234), (223, 223, 235), (218, 209, 222), (209, 193, 204), (243, 222, 230), (255, 208, 201), (214, 113, 76), (233, 89, 43), (255, 78, 41), (232, 47, 17), (227, 69, 42), (252, 93, 78), (255, 69, 74), (236, 31, 46), (237, 29, 44), (221, 23, 36), (193, 19, 28), (183, 30, 38), (195, 60, 68), (227, 81, 94), (251, 64, 84), (234, 25, 49), (241, 28, 55), (250, 38, 71), (240, 34, 79), (192, 17, 66), (112, 0, 36), (95, 0, 54), (123, 10, 101), (138, 21, 134), (110, 4, 129), (114, 4, 136), (130, 6, 139), (149, 13, 148), (179, 32, 170), (194, 55, 185), (203, 89, 201), (224, 151, 232), (252, 233, 255), (219, 224, 255), (126, 126, 190), (84, 80, 157), (172, 168, 237), (199, 196, 251), (202, 201, 235), (216, 216, 242), (227, 226, 255), (207, 206, 238), (199, 199, 227), (221, 222, 242), (221, 224, 231), (221, 224, 230), (240, 242, 255), (232, 234, 249), (237, 239, 251), (237, 240, 249), (237, 239, 250), (237, 239, 251), (237, 239, 251), (238, 239, 250), (238, 239, 248), (239, 240, 246), (0, 0, 3), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 0), (2, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 2), (0, 1, 7), (201, 212, 223), (201, 213, 227), (198, 208, 224), (197, 206, 221), (209, 213, 227), (215, 214, 226), (197, 191, 200), (178, 159, 163), (212, 171, 167), (237, 183, 174), (240, 182, 170), (235, 172, 157), (233, 166, 149), (246, 180, 165), (226, 168, 156), (235, 188, 180), (231, 198, 192), (227, 204, 204), (227, 210, 217), (238, 225, 236), (225, 211, 226), (234, 220, 236), (228, 216, 230), (242, 206, 207), (243, 156, 129), (219, 89, 48), (236, 67, 27), (220, 43, 6), (220, 67, 34), (255, 119, 100), (255, 74, 77), (225, 19, 33), (229, 11, 27), (228, 13, 30), (206, 9, 28), (202, 26, 47), (172, 18, 42), (175, 16, 45), (232, 38, 74), (226, 14, 54), (241, 31, 68), (228, 19, 60), (225, 18, 70), (215, 35, 90), (131, 3, 53), (124, 20, 81), (117, 9, 96), (112, 8, 112), (104, 10, 123), (82, 0, 104), (106, 0, 113), (129, 4, 125), (146, 5, 134), (161, 24, 150), (215, 99, 214), (235, 155, 246), (235, 205, 255), (191, 183, 235), (138, 122, 206), (138, 118, 213), (167, 149, 234), (167, 152, 220), (193, 183, 228), (216, 208, 245), (179, 171, 212), (198, 191, 232), (167, 163, 196), (195, 193, 216), (235, 236, 245), (234, 237, 244), (226, 229, 245), (239, 242, 255), (237, 239, 252), (238, 239, 249), (238, 239, 250), (238, 239, 251), (238, 239, 251), (238, 239, 250), (238, 239, 248), (239, 240, 246), (0, 0, 3), (0, 0, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 3), (0, 0, 2), (3, 0, 0), (4, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 0), (0, 2, 5), (196, 210, 221), (199, 215, 229), (190, 201, 214), (203, 208, 221), (211, 209, 221), (214, 202, 213), (219, 197, 203), (194, 150, 147), (204, 127, 109), (232, 141, 114), (228, 143, 111), (235, 156, 119), (241, 168, 127), (245, 174, 137), (255, 185, 159), (247, 179, 159), (232, 166, 148), (245, 187, 175), (241, 196, 193), (232, 200, 203), (232, 214, 218), (220, 210, 217), (226, 220, 231), (244, 219, 223), (255, 192, 177), (255, 149, 117), (247, 99, 53), (222, 59, 8), (209, 58, 13), (255, 114, 81), (255, 121, 107), (240, 62, 62), (223, 14, 27), (216, 0, 20), (207, 3, 30), (208, 25, 54), (156, 6, 31), (156, 5, 33), (205, 20, 58), (217, 13, 54), (217, 10, 46), (213, 10, 47), (201, 13, 57), (175, 16, 65), (120, 4, 57), (91, 0, 63), (105, 17, 100), (145, 58, 152), (137, 47, 146), (132, 39, 139), (91, 0, 92), (101, 0, 97), (115, 0, 106), (133, 10, 125), (171, 46, 167), (245, 143, 254), (194, 142, 226), (149, 117, 198), (168, 124, 228), (163, 116, 226), (172, 129, 228), (190, 154, 236), (212, 184, 245), (193, 171, 221), (185, 165, 215), (184, 168, 212), (201, 190, 223), (239, 234, 255), (231, 231, 241), (221, 225, 233), (215, 223, 238), (231, 238, 255), (237, 241, 253), (239, 240, 250), (239, 240, 251), (238, 239, 251), (238, 239, 251), (238, 239, 250), (238, 238, 247), (238, 238, 245), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 4), (0, 0, 3), (3, 0, 0), (4, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 0), (0, 2, 4), (195, 212, 222), (199, 217, 231), (189, 201, 214), (206, 210, 222), (213, 208, 220), (218, 203, 213), (234, 206, 211), (210, 159, 154), (220, 135, 113), (253, 154, 120), (241, 151, 107), (229, 146, 93), (240, 161, 101), (246, 166, 107), (248, 159, 112), (255, 163, 123), (255, 160, 122), (255, 174, 143), (255, 183, 161), (250, 191, 176), (247, 208, 195), (239, 211, 202), (237, 212, 209), (246, 210, 204), (255, 206, 189), (255, 182, 149), (255, 135, 83), (231, 88, 29), (226, 88, 33), (255, 125, 80), (255, 127, 100), (255, 111, 102), (231, 38, 49), (230, 20, 46), (219, 13, 50), (185, 2, 40), (142, 0, 29), (140, 4, 34), (163, 0, 36), (193, 11, 51), (193, 2, 42), (181, 0, 35), (185, 13, 60), (174, 28, 81), (102, 0, 51), (137, 50, 117), (147, 67, 146), (165, 82, 170), (204, 111, 203), (161, 64, 158), (112, 18, 107), (141, 45, 137), (123, 17, 119), (121, 4, 118), (167, 36, 166), (209, 94, 221), (173, 102, 207), (181, 126, 228), (177, 111, 228), (153, 85, 205), (158, 99, 207), (200, 151, 243), (203, 164, 237), (203, 172, 232), (202, 174, 230), (225, 203, 249), (226, 212, 245), (221, 214, 236), (234, 232, 244), (241, 244, 253), (232, 240, 254), (233, 241, 255), (236, 240, 251), (238, 239, 249), (239, 239, 250), (239, 239, 251), (239, 239, 251), (239, 239, 250), (239, 239, 248), (239, 239, 246), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 4), (0, 0, 3), (3, 0, 0), (3, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 2, 4), (197, 214, 224), (193, 212, 226), (201, 213, 226), (203, 208, 221), (211, 209, 222), (224, 212, 223), (228, 204, 210), (241, 200, 197), (250, 184, 169), (250, 172, 142), (242, 167, 119), (239, 164, 100), (244, 162, 88), (240, 146, 67), (232, 117, 43), (234, 105, 35), (238, 99, 34), (242, 108, 50), (240, 126, 75), (250, 154, 112), (255, 185, 150), (255, 198, 168), (254, 185, 158), (250, 182, 153), (249, 183, 150), (255, 191, 149), (255, 173, 117), (224, 107, 44), (229, 117, 54), (252, 141, 88), (255, 149, 115), (250, 116, 104), (254, 84, 94), (236, 44, 73), (243, 45, 88), (214, 35, 82), (144, 12, 52), (109, 0, 28), (118, 0, 21), (136, 0, 28), (161, 1, 47), (164, 0, 53), (186, 28, 88), (194, 55, 119), (148, 40, 106), (205, 115, 186), (188, 102, 181), (197, 107, 193), (200, 98, 190), (143, 36, 131), (141, 37, 133), (141, 36, 138), (125, 14, 127), (128, 8, 134), (157, 26, 167), (136, 15, 154), (147, 59, 179), (214, 138, 253), (169, 84, 209), (155, 74, 197), (183, 116, 228), (165, 111, 209), (198, 155, 236), (201, 166, 234), (202, 171, 230), (215, 192, 238), (232, 220, 252), (234, 228, 249), (244, 240, 254), (232, 230, 242), (233, 235, 249), (237, 240, 254), (236, 238, 249), (237, 238, 248), (237, 238, 249), (238, 238, 250), (239, 239, 251), (239, 239, 250), (239, 239, 248), (239, 239, 246), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 4), (0, 0, 2), (2, 0, 0), (3, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 4), (194, 209, 221), (192, 211, 225), (206, 219, 233), (203, 211, 224), (209, 210, 223), (201, 194, 205), (179, 161, 167), (206, 173, 172), (232, 180, 168), (241, 178, 153), (242, 178, 135), (239, 170, 112), (245, 165, 96), (254, 158, 81), (243, 127, 44), (220, 86, 4), (228, 80, 5), (220, 72, 0), (211, 77, 7), (217, 96, 31), (223, 114, 58), (232, 126, 76), (224, 113, 66), (225, 119, 75), (235, 143, 103), (234, 139, 98), (247, 132, 84), (249, 128, 75), (229, 117, 61), (255, 149, 101), (246, 138, 108), (244, 118, 110), (254, 91, 108), (209, 23, 60), (207, 13, 64), (218, 41, 96), (160, 22, 73), (94, 0, 21), (113, 4, 33), (119, 4, 36), (140, 10, 58), (159, 21, 81), (201, 62, 129), (230, 103, 175), (225, 122, 195), (241, 152, 229), (215, 129, 212), (215, 126, 215), (186, 86, 181), (140, 37, 137), (152, 54, 156), (96, 0, 108), (85, 0, 104), (105, 3, 131), (142, 33, 171), (184, 83, 220), (177, 99, 222), (148, 74, 195), (138, 52, 179), (152, 64, 191), (152, 74, 193), (107, 40, 146), (164, 108, 198), (183, 138, 213), (194, 160, 220), (213, 191, 236), (238, 230, 255), (239, 237, 255), (243, 242, 255), (234, 232, 244), (238, 236, 248), (237, 237, 248), (237, 238, 248), (236, 238, 248), (237, 238, 249), (237, 238, 250), (238, 239, 251), (238, 239, 250), (239, 239, 248), (240, 240, 247), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 1, 3), (0, 1, 2), (2, 0, 0), (3, 0, 0), (1, 0, 0), (0, 0, 1), (1, 0, 0), (0, 1, 5), (197, 212, 225), (198, 216, 231), (190, 204, 217), (202, 211, 224), (208, 213, 227), (199, 197, 209), (204, 193, 199), (210, 185, 184), (219, 177, 166), (248, 194, 174), (244, 185, 156), (241, 176, 139), (248, 175, 131), (249, 166, 110), (251, 155, 85), (251, 140, 65), (253, 125, 54), (241, 105, 31), (229, 93, 10), (226, 90, 6), (218, 82, 6), (223, 82, 13), (223, 73, 10), (236, 88, 34), (224, 90, 48), (234, 97, 64), (234, 77, 51), (216, 59, 32), (207, 67, 33), (255, 131, 100), (255, 140, 124), (255, 155, 160), (255, 107, 138), (229, 40, 89), (185, 0, 54), (204, 24, 87), (197, 38, 102), (119, 0, 38), (108, 2, 33), (109, 14, 43), (102, 2, 48), (132, 25, 85), (200, 84, 155), (247, 135, 213), (238, 143, 225), (221, 137, 223), (226, 147, 238), (202, 122, 219), (156, 69, 173), (184, 98, 206), (203, 125, 236), (167, 96, 209), (139, 71, 188), (134, 69, 188), (124, 60, 181), (179, 124, 244), (104, 63, 181), (81, 34, 154), (99, 27, 154), (124, 36, 166), (138, 46, 172), (163, 74, 191), (180, 104, 204), (186, 127, 208), (199, 161, 220), (230, 211, 251), (230, 229, 253), (216, 222, 237), (229, 234, 246), (236, 237, 247), (233, 231, 241), (238, 235, 245), (237, 238, 247), (236, 239, 248), (236, 238, 249), (238, 239, 251), (238, 239, 251), (238, 239, 250), (238, 239, 248), (239, 240, 246), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 1, 2), (0, 1, 1), (2, 0, 0), (3, 0, 0), (1, 0, 0), (0, 0, 1), (1, 0, 0), (0, 0, 5), (197, 211, 224), (192, 209, 225), (198, 212, 225), (207, 218, 230), (198, 207, 221), (204, 208, 220), (218, 213, 220), (202, 186, 187), (208, 177, 169), (229, 187, 175), (240, 189, 177), (255, 204, 188), (255, 194, 171), (231, 165, 129), (234, 162, 106), (240, 157, 91), (255, 155, 90), (251, 136, 62), (247, 124, 30), (250, 118, 17), (251, 111, 15), (255, 105, 18), (255, 94, 20), (255, 94, 38), (236, 80, 47), (248, 89, 73), (252, 80, 74), (189, 19, 12), (237, 83, 66), (255, 124, 107), (229, 99, 91), (255, 116, 126), (255, 89, 123), (229, 43, 92), (181, 5, 59), (176, 11, 69), (190, 36, 99), (137, 4, 60), (101, 0, 37), (97, 12, 45), (70, 0, 31), (118, 27, 86), (187, 81, 155), (229, 121, 206), (209, 110, 201), (191, 100, 197), (211, 126, 228), (176, 93, 201), (158, 75, 190), (175, 97, 216), (158, 90, 211), (160, 100, 221), (159, 107, 226), (179, 135, 250), (175, 142, 249), (130, 110, 216), (117, 112, 222), (109, 96, 213), (76, 32, 157), (88, 20, 148), (135, 49, 176), (169, 80, 197), (189, 112, 210), (192, 134, 211), (216, 183, 236), (233, 220, 255), (234, 236, 255), (230, 238, 252), (231, 238, 249), (238, 241, 250), (238, 237, 244), (243, 242, 249), (237, 238, 247), (236, 239, 248), (236, 238, 249), (236, 238, 250), (237, 239, 251), (238, 239, 250), (238, 239, 248), (239, 240, 246), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 1), (0, 2, 2), (0, 2, 0), (1, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 1), (1, 0, 0), (0, 0, 5), (202, 216, 228), (190, 208, 222), (204, 219, 232), (197, 211, 223), (188, 200, 214), (205, 213, 226), (215, 216, 225), (217, 209, 213), (220, 202, 200), (224, 195, 195), (238, 197, 203), (250, 204, 209), (243, 198, 195), (244, 200, 182), (253, 209, 171), (248, 197, 145), (251, 183, 126), (251, 168, 93), (244, 147, 44), (239, 129, 13), (244, 122, 5), (249, 115, 10), (253, 105, 25), (242, 86, 36), (216, 57, 43), (250, 91, 96), (227, 66, 77), (241, 81, 90), (255, 118, 114), (219, 66, 59), (232, 82, 77), (255, 101, 108), (244, 63, 89), (205, 27, 63), (167, 15, 52), (142, 8, 49), (141, 15, 64), (118, 4, 56), (99, 3, 51), (94, 7, 54), (89, 4, 53), (122, 30, 88), (161, 52, 128), (190, 74, 164), (183, 69, 171), (177, 68, 178), (177, 74, 190), (152, 55, 177), (123, 34, 162), (115, 35, 167), (103, 32, 167), (104, 42, 175), (96, 43, 169), (120, 81, 196), (147, 128, 227), (93, 96, 191), (90, 118, 220), (102, 128, 239), (100, 98, 218), (82, 51, 174), (171, 110, 232), (197, 126, 236), (195, 134, 220), (212, 170, 232), (214, 198, 236), (224, 223, 247), (238, 240, 255), (238, 241, 255), (226, 230, 242), (235, 238, 247), (239, 241, 247), (230, 232, 237), (235, 237, 245), (235, 238, 247), (235, 237, 248), (235, 237, 249), (236, 238, 250), (238, 239, 250), (238, 239, 248), (239, 240, 246), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 2, 1), (0, 2, 0), (1, 0, 0), (2, 0, 0), (0, 0, 0), (0, 0, 2), (1, 0, 1), (0, 0, 5), (197, 211, 223), (197, 215, 229), (193, 208, 221), (197, 211, 223), (202, 217, 231), (200, 212, 226), (204, 209, 220), (213, 212, 217), (222, 215, 211), (223, 207, 203), (231, 203, 208), (239, 207, 213), (246, 215, 215), (244, 216, 206), (238, 212, 189), (245, 215, 180), (248, 205, 161), (255, 201, 137), (252, 181, 85), (234, 148, 36), (231, 128, 14), (235, 114, 16), (249, 107, 42), (236, 80, 50), (210, 46, 53), (219, 55, 80), (241, 85, 107), (236, 82, 98), (255, 108, 111), (231, 67, 65), (241, 67, 66), (218, 40, 45), (201, 24, 42), (157, 0, 22), (125, 0, 23), (109, 4, 33), (104, 8, 44), (90, 1, 45), (86, 3, 55), (85, 7, 60), (118, 43, 92), (101, 19, 74), (115, 16, 89), (138, 30, 117), (150, 38, 138), (157, 45, 155), (141, 35, 151), (123, 25, 147), (103, 18, 146), (106, 30, 163), (105, 35, 174), (109, 45, 183), (124, 65, 197), (170, 127, 246), (144, 127, 226), (117, 131, 223), (96, 145, 245), (41, 99, 206), (82, 122, 236), (72, 82, 199), (124, 93, 207), (168, 120, 219), (209, 168, 238), (236, 210, 255), (232, 229, 255), (230, 237, 254), (232, 233, 251), (232, 232, 249), (236, 238, 251), (234, 238, 247), (231, 236, 241), (234, 239, 244), (233, 236, 244), (233, 236, 245), (234, 237, 247), (235, 237, 249), (236, 238, 250), (236, 238, 249), (238, 239, 248), (238, 240, 246), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 1), (0, 1, 0), (1, 0, 0), (2, 0, 0), (0, 0, 1), (0, 0, 2), (1, 0, 1), (0, 0, 5), (198, 210, 223), (195, 212, 227), (199, 214, 227), (199, 214, 226), (197, 213, 228), (199, 212, 227), (204, 213, 225), (209, 214, 216), (208, 211, 195), (219, 216, 194), (221, 209, 194), (225, 208, 196), (234, 217, 204), (239, 221, 210), (236, 219, 210), (238, 217, 204), (244, 215, 190), (236, 200, 155), (228, 183, 108), (236, 175, 86), (230, 147, 58), (239, 129, 59), (222, 80, 51), (212, 49, 53), (198, 25, 57), (175, 4, 44), (222, 66, 94), (255, 113, 128), (255, 120, 122), (216, 42, 41), (222, 23, 25), (208, 12, 17), (177, 12, 23), (124, 0, 6), (98, 0, 16), (84, 8, 27), (64, 0, 20), (56, 0, 27), (62, 2, 49), (65, 7, 59), (72, 19, 64), (78, 20, 69), (86, 13, 76), (99, 14, 90), (122, 28, 115), (131, 34, 130), (121, 26, 128), (106, 19, 127), (94, 21, 136), (95, 29, 153), (103, 37, 171), (119, 51, 190), (150, 80, 219), (164, 107, 236), (168, 140, 251), (133, 144, 245), (69, 129, 228), (22, 104, 206), (44, 123, 232), (58, 112, 221), (55, 60, 164), (73, 54, 138), (198, 178, 230), (230, 220, 248), (227, 236, 251), (226, 239, 250), (237, 237, 254), (239, 236, 253), (233, 237, 248), (232, 239, 247), (233, 241, 246), (232, 238, 244), (233, 238, 245), (234, 238, 247), (236, 240, 250), (236, 240, 251), (237, 239, 251), (236, 238, 249), (236, 239, 247), (237, 239, 245), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 1), (0, 1, 0), (1, 0, 0), (2, 0, 0), (0, 0, 2), (0, 0, 3), (1, 0, 1), (0, 0, 5), (198, 210, 222), (196, 212, 227), (198, 213, 225), (199, 214, 226), (198, 214, 229), (200, 215, 230), (204, 215, 228), (210, 216, 218), (205, 206, 190), (190, 186, 160), (214, 205, 180), (217, 207, 182), (226, 216, 192), (217, 205, 188), (222, 206, 201), (243, 220, 214), (246, 215, 194), (255, 222, 180), (255, 211, 145), (255, 195, 118), (248, 161, 88), (252, 136, 85), (218, 68, 60), (201, 33, 55), (185, 14, 53), (173, 5, 45), (204, 46, 70), (255, 129, 139), (248, 93, 90), (208, 37, 30), (223, 21, 20), (207, 9, 14), (154, 0, 6), (123, 1, 16), (89, 2, 21), (63, 0, 19), (54, 5, 20), (45, 0, 23), (46, 0, 37), (63, 11, 60), (71, 23, 66), (64, 12, 59), (67, 5, 62), (82, 10, 77), (100, 19, 95), (109, 24, 108), (106, 22, 111), (91, 17, 112), (77, 21, 122), (69, 19, 130), (90, 37, 161), (124, 65, 198), (129, 64, 200), (140, 86, 217), (152, 129, 244), (72, 88, 193), (12, 76, 176), (27, 119, 220), (30, 134, 239), (20, 103, 206), (25, 57, 151), (57, 59, 133), (168, 163, 203), (189, 189, 207), (217, 231, 241), (220, 234, 244), (233, 234, 251), (236, 235, 252), (229, 236, 246), (228, 239, 245), (231, 240, 247), (230, 237, 245), (233, 239, 247), (234, 238, 247), (235, 239, 249), (236, 240, 251), (236, 239, 250), (236, 239, 249), (236, 239, 247), (237, 239, 245), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 1, 0), (1, 0, 0), (2, 0, 0), (0, 0, 3), (0, 0, 4), (1, 0, 1), (0, 0, 5), (200, 213, 224), (196, 213, 226), (197, 212, 223), (198, 213, 225), (198, 214, 229), (198, 214, 229), (201, 213, 226), (208, 210, 216), (215, 202, 196), (224, 205, 189), (213, 196, 171), (227, 213, 183), (220, 211, 178), (211, 199, 173), (229, 207, 196), (244, 209, 196), (244, 191, 157), (230, 163, 110), (244, 163, 93), (255, 162, 87), (247, 132, 66), (254, 117, 74), (250, 86, 85), (194, 24, 45), (167, 10, 38), (147, 0, 18), (165, 5, 17), (255, 101, 100), (237, 88, 75), (230, 74, 58), (255, 75, 66), (210, 28, 31), (158, 0, 17), (133, 6, 33), (96, 4, 35), (65, 0, 28), (55, 9, 26), (44, 2, 21), (45, 0, 26), (66, 6, 50), (70, 10, 54), (62, 0, 48), (69, 2, 56), (85, 12, 74), (92, 15, 83), (92, 16, 89), (85, 14, 91), (70, 11, 93), (59, 21, 108), (59, 30, 126), (69, 37, 146), (85, 49, 167), (120, 75, 201), (118, 85, 209), (86, 83, 196), (57, 86, 191), (29, 89, 192), (1, 89, 190), (27, 139, 241), (36, 134, 232), (46, 93, 180), (117, 133, 199), (206, 209, 243), (227, 228, 245), (215, 228, 238), (219, 232, 243), (232, 235, 253), (234, 237, 254), (225, 238, 246), (225, 240, 245), (231, 240, 249), (232, 237, 248), (235, 239, 248), (235, 239, 248), (235, 239, 249), (235, 239, 250), (235, 239, 250), (235, 239, 249), (236, 239, 247), (237, 239, 245), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 1), (1, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 1, 0), (1, 0, 0), (2, 0, 0), (0, 0, 3), (0, 0, 4), (0, 0, 1), (0, 1, 4), (200, 213, 223), (196, 213, 225), (198, 212, 222), (199, 213, 224), (198, 214, 229), (200, 215, 230), (202, 213, 227), (209, 210, 219), (217, 203, 201), (236, 215, 203), (221, 202, 179), (222, 205, 176), (220, 207, 173), (239, 223, 193), (237, 210, 193), (255, 216, 196), (245, 184, 145), (213, 135, 78), (198, 104, 32), (202, 92, 17), (227, 99, 34), (216, 67, 25), (252, 78, 75), (228, 51, 68), (184, 25, 45), (162, 11, 26), (173, 20, 22), (255, 104, 95), (255, 124, 105), (255, 109, 88), (255, 98, 84), (210, 31, 29), (196, 32, 49), (143, 6, 35), (99, 0, 34), (73, 4, 35), (53, 5, 25), (50, 7, 27), (64, 7, 41), (76, 12, 53), (76, 11, 54), (76, 9, 55), (79, 9, 61), (82, 12, 67), (81, 13, 72), (77, 12, 77), (70, 13, 82), (59, 16, 89), (44, 20, 98), (50, 36, 122), (61, 47, 143), (66, 47, 153), (101, 75, 190), (90, 75, 191), (33, 45, 154), (25, 61, 165), (19, 72, 177), (3, 79, 183), (5, 110, 210), (59, 157, 250), (128, 183, 255), (177, 204, 255), (200, 210, 245), (214, 220, 239), (204, 217, 232), (209, 221, 236), (222, 226, 246), (224, 228, 246), (217, 231, 240), (220, 235, 241), (230, 236, 248), (234, 236, 249), (235, 239, 249), (235, 239, 248), (234, 238, 248), (234, 238, 249), (235, 239, 250), (235, 239, 249), (236, 239, 247), (237, 239, 245), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 1), (1, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 3), (0, 0, 4), (0, 0, 1), (0, 1, 4), (198, 211, 219), (195, 212, 222), (199, 212, 221), (201, 214, 224), (201, 216, 230), (202, 216, 232), (205, 215, 230), (209, 213, 222), (219, 216, 211), (223, 213, 199), (225, 209, 192), (221, 202, 180), (230, 210, 184), (237, 213, 187), (243, 212, 191), (255, 214, 187), (254, 198, 158), (234, 163, 108), (239, 154, 81), (240, 136, 58), (250, 123, 53), (199, 47, 0), (203, 23, 8), (203, 14, 20), (201, 25, 38), (172, 12, 21), (156, 17, 11), (209, 72, 56), (253, 99, 79), (252, 81, 61), (255, 81, 65), (255, 68, 62), (213, 36, 46), (149, 0, 20), (104, 0, 24), (80, 2, 32), (55, 1, 26), (57, 8, 36), (74, 14, 51), (75, 10, 51), (80, 13, 55), (88, 21, 64), (86, 17, 64), (77, 11, 60), (72, 13, 67), (64, 14, 73), (53, 12, 78), (46, 17, 88), (31, 17, 93), (46, 41, 122), (46, 43, 130), (45, 41, 135), (54, 46, 148), (45, 46, 151), (14, 36, 139), (0, 28, 132), (0, 36, 146), (4, 61, 169), (25, 108, 209), (54, 136, 227), (95, 150, 227), (161, 195, 255), (185, 205, 246), (186, 200, 229), (194, 209, 233), (200, 212, 234), (212, 217, 240), (218, 222, 241), (216, 227, 238), (224, 234, 243), (236, 238, 252), (240, 239, 254), (235, 239, 249), (233, 239, 247), (234, 238, 248), (234, 238, 249), (234, 238, 249), (235, 239, 249), (236, 239, 247), (237, 239, 245), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 1), (1, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 3), (0, 0, 4), (0, 0, 1), (0, 1, 4), (198, 212, 220), (196, 213, 222), (199, 212, 220), (201, 212, 223), (199, 212, 227), (199, 212, 229), (202, 211, 227), (205, 209, 219), (201, 201, 199), (205, 199, 191), (216, 202, 192), (236, 214, 199), (240, 213, 187), (250, 214, 181), (255, 224, 187), (255, 213, 174), (255, 197, 157), (255, 174, 124), (255, 179, 110), (255, 169, 91), (255, 152, 74), (239, 92, 30), (191, 18, 0), (207, 24, 12), (196, 19, 18), (159, 0, 0), (137, 3, 0), (145, 14, 0), (216, 65, 47), (214, 46, 27), (226, 43, 26), (230, 43, 33), (216, 36, 39), (169, 13, 26), (121, 6, 26), (86, 4, 28), (62, 3, 30), (66, 11, 43), (82, 13, 52), (87, 10, 53), (91, 14, 59), (98, 19, 66), (97, 16, 65), (86, 12, 63), (74, 14, 67), (60, 14, 71), (49, 16, 80), (45, 24, 93), (44, 35, 108), (45, 44, 121), (32, 38, 117), (18, 27, 111), (17, 26, 118), (14, 32, 129), (0, 31, 129), (0, 43, 146), (0, 42, 151), (0, 50, 158), (22, 89, 187), (28, 91, 179), (81, 124, 201), (172, 199, 255), (185, 201, 253), (192, 204, 246), (193, 207, 242), (196, 210, 239), (206, 216, 240), (214, 223, 241), (217, 228, 240), (227, 234, 245), (237, 236, 251), (237, 235, 250), (232, 236, 246), (232, 238, 246), (233, 238, 248), (234, 238, 249), (234, 238, 249), (234, 238, 248), (235, 238, 246), (237, 239, 245), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 1), (1, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (2, 0, 0), (1, 0, 0), (0, 1, 3), (0, 1, 4), (0, 1, 1), (0, 1, 4), (198, 212, 220), (197, 214, 223), (200, 213, 221), (201, 212, 222), (197, 210, 225), (197, 209, 226), (199, 206, 223), (202, 205, 219), (210, 207, 215), (210, 202, 205), (230, 217, 218), (233, 212, 200), (237, 205, 171), (255, 209, 157), (241, 166, 101), (255, 162, 102), (255, 138, 99), (225, 89, 50), (245, 115, 54), (255, 149, 71), (255, 131, 41), (255, 131, 48), (241, 91, 32), (233, 74, 34), (210, 50, 24), (171, 18, 2), (151, 13, 2), (133, 0, 0), (188, 46, 33), (189, 39, 23), (195, 32, 15), (191, 20, 7), (221, 46, 43), (180, 24, 27), (127, 10, 18), (85, 0, 14), (60, 0, 23), (72, 11, 43), (104, 19, 58), (125, 28, 73), (121, 21, 74), (123, 21, 78), (138, 35, 92), (136, 43, 100), (98, 27, 84), (64, 13, 72), (55, 20, 85), (53, 32, 100), (57, 45, 117), (28, 28, 101), (28, 40, 113), (23, 45, 120), (5, 33, 115), (5, 42, 130), (0, 42, 137), (0, 60, 159), (0, 62, 164), (21, 92, 192), (68, 126, 219), (98, 138, 225), (149, 167, 249), (184, 189, 255), (194, 193, 255), (193, 194, 252), (189, 198, 245), (189, 203, 239), (195, 213, 236), (205, 223, 238), (214, 228, 239), (223, 231, 243), (228, 227, 243), (224, 222, 237), (230, 234, 244), (230, 237, 245), (233, 239, 248), (233, 238, 249), (233, 237, 248), (233, 237, 247), (235, 238, 246), (237, 239, 245), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 1), (1, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 3), (0, 1, 3), (0, 1, 1), (0, 2, 4), (197, 210, 218), (197, 212, 223), (200, 213, 222), (201, 213, 224), (199, 212, 226), (200, 212, 227), (202, 211, 227), (206, 211, 225), (211, 209, 220), (219, 212, 220), (223, 210, 220), (217, 190, 183), (255, 206, 164), (237, 161, 99), (210, 100, 32), (230, 92, 35), (218, 62, 31), (189, 28, 1), (197, 47, 1), (237, 95, 32), (226, 90, 13), (236, 100, 25), (242, 97, 40), (236, 89, 45), (232, 86, 51), (204, 61, 36), (180, 41, 28), (166, 32, 23), (149, 20, 8), (149, 20, 6), (144, 10, 0), (160, 20, 6), (176, 30, 23), (135, 1, 0), (99, 0, 0), (76, 0, 8), (56, 0, 18), (71, 6, 37), (111, 16, 56), (136, 25, 73), (135, 22, 76), (144, 29, 87), (193, 75, 135), (211, 104, 164), (144, 66, 123), (75, 23, 80), (50, 18, 77), (39, 22, 84), (29, 20, 85), (21, 23, 90), (9, 25, 93), (20, 47, 120), (11, 48, 129), (5, 53, 143), (4, 66, 164), (1, 76, 176), (8, 95, 191), (45, 124, 218), (121, 171, 255), (122, 149, 239), (138, 146, 231), (162, 162, 242), (168, 170, 246), (178, 183, 251), (181, 192, 249), (181, 198, 243), (187, 212, 241), (200, 225, 244), (215, 232, 249), (225, 234, 250), (227, 228, 246), (220, 220, 236), (227, 232, 243), (230, 237, 245), (233, 240, 249), (234, 240, 250), (232, 237, 248), (232, 236, 246), (233, 237, 245), (236, 239, 245), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (1, 0, 1), (1, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 2), (1, 0, 3), (0, 0, 2), (0, 0, 1), (0, 1, 1), (0, 1, 5), (201, 211, 221), (199, 211, 225), (199, 211, 225), (200, 214, 226), (200, 215, 227), (201, 216, 228), (203, 215, 230), (205, 214, 228), (201, 206, 212), (215, 212, 220), (214, 200, 217), (232, 194, 192), (251, 176, 127), (214, 100, 37), (202, 50, 3), (209, 37, 6), (200, 31, 15), (188, 24, 9), (177, 20, 0), (183, 29, 0), (196, 39, 0), (191, 34, 0), (194, 41, 10), (189, 43, 16), (184, 49, 19), (172, 42, 15), (198, 65, 46), (180, 52, 38), (132, 17, 5), (117, 12, 0), (103, 7, 0), (95, 2, 0), (96, 0, 0), (106, 18, 14), (78, 9, 10), (55, 0, 6), (49, 0, 14), (63, 0, 26), (108, 8, 51), (130, 13, 63), (153, 35, 84), (226, 105, 157), (195, 69, 127), (195, 83, 142), (128, 49, 104), (66, 16, 67), (45, 22, 70), (26, 19, 68), (15, 15, 67), (7, 15, 73), (13, 29, 96), (8, 35, 112), (2, 40, 130), (3, 58, 157), (0, 74, 181), (2, 90, 194), (12, 106, 197), (46, 126, 215), (93, 137, 234), (133, 156, 252), (127, 140, 228), (147, 159, 242), (146, 167, 246), (153, 176, 250), (169, 187, 255), (175, 196, 252), (185, 216, 255), (193, 224, 253), (211, 229, 255), (213, 223, 250), (223, 229, 251), (234, 239, 255), (229, 236, 246), (230, 237, 245), (231, 238, 247), (231, 238, 248), (232, 238, 248), (232, 238, 247), (234, 239, 246), (236, 240, 245), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (1, 0, 0), (1, 0, 0), (2, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (202, 210, 221), (200, 210, 225), (198, 211, 226), (198, 213, 226), (200, 216, 226), (200, 215, 226), (200, 214, 230), (201, 213, 227), (204, 213, 220), (221, 221, 229), (223, 210, 225), (243, 200, 193), (255, 172, 115), (215, 82, 16), (216, 42, 6), (216, 29, 13), (205, 33, 26), (157, 0, 0), (156, 8, 0), (158, 12, 0), (172, 20, 2), (170, 19, 0), (147, 3, 0), (141, 8, 0), (141, 23, 0), (162, 48, 2), (175, 55, 12), (174, 55, 16), (138, 28, 0), (134, 32, 3), (120, 27, 3), (97, 9, 0), (80, 0, 0), (71, 0, 0), (74, 8, 11), (66, 6, 15), (66, 5, 20), (76, 0, 26), (114, 11, 50), (177, 60, 106), (220, 101, 147), (252, 131, 181), (203, 78, 136), (165, 57, 116), (108, 35, 90), (49, 8, 58), (31, 16, 63), (19, 20, 67), (12, 19, 70), (4, 19, 76), (0, 25, 92), (2, 40, 119), (14, 66, 158), (22, 91, 193), (20, 111, 220), (28, 131, 236), (49, 156, 244), (68, 162, 248), (74, 138, 234), (96, 143, 241), (110, 154, 245), (109, 154, 239), (112, 166, 245), (116, 168, 244), (127, 166, 240), (126, 167, 232), (126, 182, 230), (151, 208, 246), (172, 215, 250), (176, 205, 236), (209, 225, 248), (201, 211, 227), (227, 237, 247), (229, 238, 245), (231, 238, 247), (231, 238, 248), (231, 238, 248), (232, 238, 247), (233, 239, 246), (234, 239, 244), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (1, 0, 0), (2, 0, 0), (2, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (202, 210, 221), (200, 210, 225), (198, 211, 226), (198, 213, 226), (199, 215, 225), (199, 214, 225), (199, 213, 229), (199, 212, 228), (205, 217, 229), (192, 196, 204), (225, 213, 216), (247, 204, 183), (248, 157, 93), (238, 104, 35), (189, 13, 0), (207, 22, 10), (192, 27, 24), (154, 8, 9), (135, 9, 9), (134, 16, 13), (140, 20, 11), (129, 10, 0), (131, 17, 0), (140, 34, 0), (207, 112, 46), (213, 121, 39), (204, 105, 20), (219, 113, 30), (217, 102, 26), (211, 90, 26), (188, 63, 17), (157, 33, 5), (138, 23, 12), (103, 0, 0), (87, 0, 2), (102, 14, 27), (106, 15, 32), (105, 9, 32), (122, 17, 48), (191, 79, 118), (247, 130, 175), (255, 140, 192), (212, 100, 157), (128, 36, 95), (76, 20, 76), (38, 9, 64), (25, 18, 73), (12, 19, 75), (15, 29, 90), (7, 33, 98), (0, 44, 115), (19, 80, 159), (33, 110, 199), (17, 109, 208), (11, 121, 226), (29, 150, 251), (42, 168, 255), (58, 180, 255), (56, 165, 255), (56, 158, 252), (54, 155, 247), (38, 137, 224), (50, 148, 227), (66, 156, 231), (91, 166, 241), (76, 153, 222), (63, 164, 219), (43, 147, 192), (74, 164, 199), (135, 202, 229), (196, 229, 250), (212, 227, 242), (226, 237, 247), (229, 238, 245), (231, 238, 247), (231, 238, 248), (231, 238, 248), (232, 238, 247), (232, 238, 245), (234, 239, 244), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (1, 0, 0), (1, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (202, 210, 221), (200, 210, 225), (198, 211, 226), (198, 213, 226), (199, 215, 225), (199, 214, 225), (199, 213, 229), (200, 213, 230), (201, 216, 230), (208, 215, 225), (225, 216, 219), (222, 183, 162), (182, 98, 37), (213, 85, 19), (225, 57, 19), (216, 35, 15), (176, 9, 0), (151, 1, 0), (134, 3, 0), (118, 0, 0), (124, 6, 0), (128, 14, 0), (157, 47, 21), (201, 98, 53), (211, 117, 44), (213, 121, 30), (227, 130, 33), (237, 131, 30), (245, 127, 27), (238, 109, 18), (235, 94, 24), (229, 85, 39), (173, 38, 17), (125, 0, 0), (111, 0, 4), (127, 14, 33), (127, 11, 35), (133, 20, 49), (102, 0, 29), (160, 55, 93), (207, 94, 140), (218, 105, 157), (213, 110, 166), (123, 42, 100), (65, 19, 74), (37, 17, 72), (23, 22, 79), (10, 22, 81), (9, 27, 90), (1, 31, 99), (0, 45, 118), (21, 87, 167), (28, 109, 199), (2, 97, 197), (0, 105, 211), (7, 129, 232), (13, 144, 234), (11, 146, 231), (19, 152, 239), (21, 152, 241), (13, 141, 233), (20, 144, 233), (17, 138, 219), (26, 139, 216), (64, 164, 240), (64, 165, 236), (39, 156, 217), (29, 146, 196), (70, 171, 206), (108, 182, 208), (168, 205, 226), (188, 204, 220), (226, 237, 247), (230, 238, 245), (231, 238, 247), (231, 238, 247), (231, 237, 247), (231, 237, 246), (233, 238, 245), (235, 239, 244), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (201, 209, 220), (199, 209, 224), (198, 211, 226), (198, 213, 226), (199, 215, 225), (200, 215, 226), (200, 214, 230), (200, 214, 231), (197, 213, 229), (211, 220, 235), (215, 210, 223), (239, 206, 200), (232, 161, 116), (179, 67, 9), (200, 48, 0), (230, 55, 15), (204, 26, 0), (189, 15, 0), (173, 8, 0), (180, 24, 10), (177, 29, 11), (161, 21, 0), (188, 57, 30), (200, 78, 38), (221, 107, 46), (220, 109, 35), (223, 109, 28), (215, 97, 6), (238, 118, 12), (255, 138, 31), (255, 128, 34), (237, 89, 16), (186, 40, 0), (153, 10, 0), (120, 0, 0), (142, 5, 31), (148, 11, 47), (136, 9, 51), (107, 3, 45), (119, 21, 64), (154, 47, 93), (159, 52, 102), (185, 88, 141), (130, 54, 108), (68, 25, 77), (38, 21, 72), (18, 21, 72), (13, 27, 82), (13, 32, 92), (3, 31, 97), (0, 34, 107), (0, 53, 136), (2, 68, 162), (0, 77, 181), (2, 95, 206), (0, 103, 212), (0, 119, 218), (11, 143, 233), (27, 165, 248), (18, 153, 237), (2, 127, 218), (7, 128, 220), (1, 124, 210), (12, 133, 214), (28, 144, 221), (37, 148, 220), (40, 148, 212), (69, 163, 216), (129, 202, 238), (151, 202, 229), (171, 200, 224), (169, 183, 202), (227, 237, 247), (230, 237, 244), (230, 237, 245), (231, 237, 246), (231, 236, 246), (232, 236, 246), (233, 237, 245), (234, 237, 243), (0, 0, 3), (0, 0, 1), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (200, 208, 219), (199, 209, 224), (199, 212, 227), (199, 214, 227), (199, 215, 225), (200, 215, 226), (201, 215, 231), (202, 216, 234), (197, 214, 231), (209, 219, 235), (217, 214, 225), (232, 207, 194), (255, 218, 162), (239, 152, 72), (209, 89, 4), (255, 115, 30), (255, 118, 38), (217, 53, 0), (220, 53, 4), (210, 44, 5), (190, 28, 0), (183, 26, 0), (174, 24, 0), (176, 33, 2), (191, 54, 12), (187, 54, 3), (192, 59, 2), (229, 100, 25), (247, 128, 24), (254, 135, 16), (255, 131, 13), (248, 110, 9), (221, 78, 10), (191, 46, 8), (187, 40, 31), (176, 28, 41), (172, 22, 51), (144, 8, 45), (104, 0, 37), (97, 6, 45), (113, 18, 60), (113, 20, 65), (134, 51, 98), (104, 39, 87), (56, 19, 64), (38, 24, 67), (19, 22, 66), (10, 22, 70), (16, 32, 85), (5, 28, 89), (0, 31, 103), (2, 43, 126), (0, 50, 146), (0, 65, 171), (6, 87, 201), (0, 99, 211), (10, 126, 227), (23, 152, 243), (7, 143, 225), (0, 119, 201), (1, 122, 213), (4, 122, 213), (2, 125, 210), (3, 127, 205), (8, 128, 199), (32, 141, 208), (83, 174, 237), (114, 186, 237), (148, 199, 234), (183, 217, 243), (207, 229, 252), (223, 236, 254), (227, 237, 247), (230, 237, 244), (230, 237, 245), (231, 237, 245), (231, 236, 246), (232, 236, 245), (233, 236, 244), (235, 237, 242), (0, 0, 3), (0, 0, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 1), (0, 0, 2), (0, 0, 2), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (200, 208, 219), (199, 209, 224), (199, 212, 227), (199, 214, 227), (199, 215, 225), (200, 215, 226), (201, 215, 231), (202, 216, 234), (199, 216, 235), (203, 214, 226), (218, 215, 210), (241, 222, 182), (252, 216, 123), (255, 211, 82), (255, 193, 45), (255, 187, 35), (255, 171, 27), (246, 124, 0), (246, 107, 11), (240, 88, 12), (221, 60, 0), (208, 42, 0), (201, 33, 4), (187, 19, 0), (176, 13, 0), (179, 21, 2), (172, 18, 0), (182, 42, 0), (211, 97, 2), (244, 140, 16), (255, 151, 11), (252, 138, 5), (233, 109, 5), (239, 106, 31), (246, 105, 60), (228, 80, 61), (192, 39, 42), (147, 8, 24), (114, 8, 27), (85, 0, 25), (83, 6, 40), (85, 15, 53), (86, 23, 62), (65, 16, 54), (40, 10, 45), (32, 18, 52), (19, 18, 52), (12, 17, 55), (6, 14, 59), (0, 12, 67), (6, 25, 93), (14, 44, 125), (13, 57, 152), (5, 65, 171), (3, 80, 195), (11, 106, 218), (25, 140, 239), (36, 163, 252), (12, 141, 225), (0, 111, 195), (0, 112, 202), (16, 130, 218), (26, 149, 226), (44, 166, 234), (44, 157, 217), (63, 158, 214), (91, 159, 214), (151, 199, 245), (181, 216, 246), (187, 211, 232), (205, 222, 240), (208, 221, 235), (227, 237, 246), (230, 238, 245), (230, 237, 245), (231, 237, 245), (231, 237, 245), (231, 235, 243), (233, 236, 243), (235, 237, 242), (0, 0, 3), (0, 0, 1), (0, 1, 0), (0, 1, 0), (0, 1, 0), (0, 0, 1), (0, 0, 2), (0, 0, 2), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (200, 208, 219), (200, 210, 225), (199, 212, 227), (199, 214, 227), (199, 215, 225), (199, 214, 225), (200, 214, 230), (201, 215, 233), (203, 219, 236), (207, 217, 218), (221, 215, 184), (242, 223, 149), (254, 223, 97), (237, 196, 35), (243, 194, 15), (248, 187, 3), (255, 181, 5), (255, 174, 15), (255, 151, 19), (250, 117, 6), (246, 97, 3), (234, 73, 1), (226, 55, 11), (214, 40, 15), (199, 29, 15), (177, 12, 0), (173, 14, 0), (167, 28, 0), (223, 117, 14), (255, 165, 27), (252, 162, 6), (255, 158, 7), (254, 144, 22), (250, 127, 33), (248, 112, 48), (229, 81, 44), (198, 39, 27), (193, 45, 48), (143, 29, 36), (102, 11, 26), (81, 2, 32), (83, 14, 51), (68, 10, 44), (53, 9, 41), (40, 13, 41), (18, 4, 31), (11, 7, 34), (16, 19, 51), (9, 16, 54), (5, 17, 66), (7, 25, 88), (10, 39, 116), (21, 63, 156), (19, 74, 180), (8, 76, 192), (16, 100, 214), (33, 138, 238), (54, 170, 255), (57, 177, 255), (25, 142, 230), (0, 92, 183), (2, 109, 196), (3, 118, 195), (38, 151, 219), (88, 190, 249), (113, 194, 246), (139, 189, 236), (176, 205, 245), (205, 225, 253), (218, 232, 252), (210, 222, 239), (223, 234, 247), (227, 237, 246), (229, 238, 245), (230, 237, 245), (230, 237, 245), (230, 236, 244), (231, 235, 243), (233, 236, 242), (234, 236, 240), (0, 0, 2), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 1, 0), (0, 1, 1), (0, 0, 3), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (201, 209, 220), (200, 210, 225), (198, 211, 226), (198, 213, 226), (199, 215, 225), (200, 215, 226), (200, 214, 230), (202, 215, 230), (202, 216, 227), (214, 220, 203), (236, 224, 158), (243, 216, 104), (249, 209, 54), (248, 199, 21), (239, 184, 4), (251, 189, 10), (255, 186, 11), (255, 177, 10), (251, 156, 2), (255, 145, 4), (255, 134, 7), (254, 112, 9), (246, 89, 18), (226, 63, 15), (204, 44, 11), (170, 16, 0), (171, 24, 0), (212, 86, 10), (254, 159, 31), (255, 177, 17), (255, 187, 18), (255, 178, 21), (251, 154, 30), (250, 138, 44), (248, 117, 51), (236, 86, 45), (236, 67, 52), (218, 56, 53), (158, 27, 27), (125, 15, 26), (124, 22, 54), (109, 21, 61), (74, 6, 40), (56, 7, 37), (32, 2, 27), (24, 9, 32), (9, 4, 28), (14, 18, 46), (2, 15, 49), (0, 16, 61), (2, 31, 89), (0, 37, 110), (7, 54, 143), (8, 61, 165), (11, 68, 184), (17, 84, 200), (20, 105, 210), (23, 121, 219), (34, 141, 236), (68, 176, 255), (39, 141, 233), (0, 90, 180), (0, 76, 163), (10, 107, 185), (75, 161, 227), (140, 206, 255), (175, 211, 253), (199, 215, 248), (210, 219, 245), (223, 228, 250), (231, 236, 255), (230, 236, 252), (231, 241, 250), (229, 239, 246), (228, 237, 245), (228, 235, 244), (231, 237, 245), (234, 238, 246), (234, 237, 243), (232, 234, 238), (0, 1, 2), (0, 1, 0), (0, 1, 0), (0, 1, 0), (0, 1, 0), (0, 1, 1), (0, 0, 3), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (201, 209, 220), (200, 210, 225), (198, 211, 226), (198, 213, 226), (199, 215, 225), (200, 215, 226), (200, 214, 230), (201, 214, 228), (208, 220, 227), (217, 220, 201), (228, 216, 150), (225, 198, 89), (229, 189, 41), (237, 186, 16), (242, 183, 9), (255, 192, 15), (255, 187, 12), (249, 170, 0), (249, 161, 0), (255, 156, 6), (255, 145, 9), (253, 120, 6), (247, 97, 12), (226, 69, 7), (203, 50, 2), (209, 61, 17), (203, 62, 10), (220, 98, 17), (255, 176, 46), (255, 194, 35), (255, 191, 25), (249, 173, 18), (254, 163, 39), (248, 140, 43), (251, 120, 48), (250, 98, 51), (253, 80, 59), (220, 50, 44), (190, 46, 43), (181, 54, 63), (171, 52, 81), (141, 37, 74), (115, 33, 64), (92, 30, 57), (52, 7, 31), (44, 15, 38), (18, 3, 27), (9, 7, 35), (4, 14, 48), (4, 26, 68), (6, 37, 92), (0, 34, 103), (0, 45, 129), (4, 52, 150), (15, 64, 173), (23, 79, 191), (15, 86, 191), (15, 100, 199), (12, 109, 204), (19, 120, 212), (71, 168, 255), (42, 136, 226), (0, 74, 167), (18, 107, 193), (56, 140, 212), (125, 190, 246), (171, 205, 243), (195, 209, 236), (195, 200, 224), (220, 222, 244), (228, 233, 254), (224, 231, 248), (221, 231, 241), (226, 236, 244), (229, 239, 248), (230, 238, 248), (230, 236, 245), (231, 235, 243), (233, 236, 242), (234, 236, 240), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 1, 0), (0, 1, 0), (0, 0, 1), (0, 0, 2), (0, 0, 2), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (201, 209, 220), (200, 210, 225), (198, 211, 226), (198, 213, 226), (199, 215, 225), (199, 214, 225), (200, 214, 230), (202, 214, 228), (207, 216, 223), (217, 220, 211), (227, 218, 186), (226, 207, 141), (234, 203, 97), (246, 202, 63), (253, 195, 32), (255, 193, 17), (255, 185, 10), (255, 166, 0), (255, 168, 18), (255, 157, 22), (252, 133, 13), (239, 106, 3), (241, 92, 8), (233, 78, 11), (218, 66, 10), (227, 79, 31), (193, 48, 3), (179, 53, 0), (233, 142, 33), (250, 180, 42), (248, 184, 34), (244, 172, 27), (249, 158, 35), (247, 135, 34), (255, 122, 42), (252, 97, 43), (251, 78, 54), (228, 56, 49), (205, 52, 48), (195, 56, 62), (157, 26, 48), (139, 22, 50), (141, 43, 68), (134, 50, 75), (108, 36, 63), (74, 18, 46), (37, 1, 29), (23, 7, 37), (14, 16, 50), (11, 26, 68), (5, 26, 80), (2, 31, 97), (13, 50, 127), (12, 55, 141), (15, 60, 154), (11, 63, 162), (8, 72, 171), (16, 92, 188), (12, 101, 192), (15, 111, 197), (16, 111, 194), (12, 106, 192), (6, 97, 193), (20, 111, 203), (10, 103, 179), (81, 159, 216), (155, 201, 235), (180, 202, 225), (208, 214, 236), (207, 209, 230), (216, 226, 245), (229, 242, 255), (228, 241, 251), (228, 240, 248), (228, 238, 248), (227, 236, 246), (229, 236, 246), (232, 238, 246), (233, 236, 243), (233, 235, 239), (0, 1, 1), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 2), (0, 0, 2), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (201, 209, 220), (199, 209, 224), (198, 211, 226), (198, 213, 226), (199, 215, 225), (199, 214, 225), (200, 214, 230), (202, 214, 229), (203, 213, 222), (210, 216, 217), (219, 217, 209), (230, 217, 183), (244, 217, 140), (252, 208, 94), (251, 187, 39), (249, 167, 5), (255, 168, 11), (252, 146, 0), (251, 143, 11), (238, 125, 6), (234, 113, 5), (229, 97, 3), (225, 79, 1), (216, 63, 0), (218, 65, 11), (193, 41, 0), (173, 22, 0), (168, 37, 0), (213, 119, 23), (254, 183, 58), (255, 209, 67), (255, 192, 52), (248, 155, 32), (248, 132, 29), (254, 116, 35), (238, 83, 29), (228, 62, 38), (231, 65, 57), (218, 65, 58), (212, 71, 70), (159, 27, 40), (118, 0, 16), (156, 47, 66), (180, 81, 102), (154, 63, 89), (105, 31, 58), (80, 33, 60), (33, 10, 39), (11, 12, 44), (10, 25, 64), (7, 26, 77), (15, 39, 100), (21, 52, 123), (7, 46, 123), (9, 53, 136), (13, 64, 152), (8, 69, 159), (4, 76, 166), (13, 96, 183), (7, 98, 181), (0, 81, 160), (1, 99, 180), (0, 93, 182), (0, 92, 178), (0, 99, 171), (61, 152, 207), (154, 217, 252), (171, 211, 236), (192, 215, 238), (201, 216, 237), (221, 237, 254), (211, 227, 241), (215, 229, 239), (221, 234, 243), (227, 238, 248), (227, 237, 247), (228, 235, 245), (228, 234, 242), (231, 235, 242), (234, 236, 240), (0, 1, 1), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (201, 209, 220), (199, 209, 224), (198, 211, 226), (198, 213, 226), (198, 214, 224), (199, 214, 225), (200, 214, 230), (200, 214, 230), (203, 220, 232), (202, 216, 225), (206, 213, 219), (224, 217, 200), (242, 215, 155), (249, 198, 101), (252, 173, 46), (250, 148, 12), (248, 131, 8), (241, 117, 4), (231, 108, 3), (210, 88, 0), (215, 90, 0), (220, 88, 2), (213, 70, 1), (203, 52, 0), (202, 45, 2), (182, 22, 0), (171, 13, 0), (171, 33, 0), (239, 138, 49), (255, 202, 80), (255, 195, 53), (247, 176, 34), (251, 154, 30), (244, 124, 22), (236, 96, 21), (212, 60, 13), (193, 39, 21), (191, 39, 33), (228, 85, 70), (244, 110, 98), (210, 85, 87), (148, 31, 41), (163, 50, 63), (174, 66, 83), (160, 56, 79), (125, 41, 66), (82, 31, 54), (31, 12, 35), (13, 22, 47), (9, 31, 64), (5, 26, 71), (15, 37, 93), (16, 44, 109), (5, 41, 112), (7, 52, 127), (14, 68, 146), (10, 76, 154), (0, 73, 153), (2, 78, 163), (0, 73, 156), (0, 88, 165), (1, 108, 180), (27, 131, 202), (18, 123, 189), (47, 156, 213), (89, 192, 241), (120, 206, 247), (135, 205, 239), (152, 206, 234), (182, 220, 242), (197, 220, 234), (219, 234, 244), (225, 239, 249), (224, 238, 248), (223, 236, 246), (223, 234, 244), (226, 234, 244), (231, 237, 245), (232, 236, 243), (233, 235, 239), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 1, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (201, 209, 220), (199, 209, 224), (198, 211, 226), (198, 213, 226), (198, 214, 224), (199, 214, 225), (200, 214, 230), (200, 215, 230), (201, 219, 231), (201, 218, 229), (205, 216, 228), (223, 220, 211), (235, 211, 158), (237, 187, 98), (242, 161, 43), (240, 135, 10), (241, 119, 10), (241, 111, 13), (229, 100, 6), (210, 81, 0), (205, 75, 0), (216, 82, 1), (216, 76, 8), (212, 64, 11), (195, 40, 2), (190, 31, 6), (172, 15, 0), (157, 17, 0), (226, 116, 44), (255, 174, 71), (245, 168, 44), (250, 170, 39), (255, 155, 33), (254, 134, 29), (234, 99, 17), (209, 65, 12), (185, 41, 21), (158, 18, 10), (221, 88, 73), (226, 101, 89), (163, 46, 46), (139, 26, 35), (148, 36, 48), (153, 42, 59), (168, 56, 79), (163, 67, 93), (81, 20, 44), (47, 20, 43), (21, 27, 51), (11, 33, 64), (7, 28, 72), (11, 36, 91), (9, 42, 104), (8, 49, 118), (8, 59, 132), (7, 69, 143), (6, 81, 155), (6, 88, 163), (6, 87, 167), (14, 104, 183), (6, 114, 186), (24, 139, 204), (91, 201, 255), (84, 197, 249), (70, 192, 238), (56, 177, 221), (65, 178, 222), (102, 201, 242), (121, 201, 234), (150, 210, 234), (185, 221, 236), (210, 232, 243), (220, 237, 248), (223, 237, 248), (224, 237, 247), (225, 236, 246), (228, 236, 246), (231, 237, 245), (232, 237, 243), (233, 235, 239), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 1), (0, 0, 1), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 4), (1, 0, 4), (0, 0, 1), (0, 0, 0), (0, 1, 1), (0, 1, 5), (201, 209, 220), (199, 209, 224), (198, 211, 226), (197, 212, 225), (198, 214, 224), (199, 214, 225), (200, 214, 230), (200, 215, 229), (198, 214, 223), (201, 216, 223), (204, 216, 223), (218, 219, 206), (226, 208, 152), (224, 183, 91), (224, 156, 33), (214, 123, 0), (224, 115, 0), (219, 98, 0), (212, 85, 0), (218, 86, 0), (207, 71, 0), (219, 81, 1), (221, 81, 6), (208, 65, 4), (187, 41, 1), (154, 6, 0), (152, 7, 0), (156, 19, 2), (188, 64, 20), (221, 109, 41), (249, 147, 57), (248, 148, 43), (254, 150, 34), (255, 150, 35), (251, 128, 26), (232, 101, 26), (196, 62, 28), (165, 33, 22), (193, 69, 61), (173, 56, 55), (144, 34, 43), (127, 21, 35), (139, 33, 50), (146, 36, 57), (152, 33, 62), (164, 56, 88), (119, 41, 71), (67, 22, 51), (25, 16, 45), (15, 28, 63), (21, 42, 88), (21, 52, 108), (2, 46, 110), (1, 55, 126), (5, 70, 145), (13, 89, 166), (21, 110, 188), (17, 113, 190), (23, 118, 193), (27, 128, 199), (25, 142, 206), (41, 163, 219), (48, 164, 213), (48, 171, 213), (24, 165, 202), (21, 169, 208), (29, 170, 216), (58, 185, 230), (107, 209, 246), (132, 211, 240), (163, 218, 238), (177, 213, 227), (176, 198, 210), (200, 215, 226), (223, 236, 247), (230, 241, 252), (227, 236, 245), (224, 231, 239), (229, 234, 240), (235, 237, 241), (0, 0, 0), (0, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 3), (0, 0, 3), (0, 0, 1), (0, 0, 0), (0, 1, 0), (0, 1, 5), (201, 209, 220), (198, 210, 224), (198, 211, 227), (197, 212, 226), (198, 213, 224), (199, 214, 225), (200, 215, 229), (200, 215, 228), (201, 217, 225), (202, 217, 222), (201, 213, 219), (214, 217, 208), (224, 214, 171), (231, 201, 125), (237, 182, 73), (225, 150, 22), (213, 122, 0), (217, 112, 0), (232, 120, 3), (255, 141, 36), (238, 108, 15), (243, 108, 24), (254, 117, 37), (243, 105, 40), (219, 78, 41), (164, 23, 4), (141, 1, 0), (183, 44, 32), (239, 100, 75), (234, 99, 60), (224, 96, 44), (202, 81, 10), (234, 121, 25), (239, 128, 21), (244, 126, 26), (235, 113, 37), (180, 55, 22), (163, 40, 33), (149, 35, 37), (133, 26, 35), (135, 32, 46), (130, 27, 45), (141, 32, 52), (155, 38, 62), (174, 47, 76), (164, 46, 77), (150, 60, 89), (75, 19, 48), (36, 20, 51), (11, 19, 57), (19, 37, 86), (25, 56, 113), (7, 56, 118), (6, 68, 135), (10, 81, 153), (23, 103, 179), (36, 127, 206), (32, 131, 208), (37, 138, 209), (29, 137, 201), (32, 151, 207), (35, 154, 202), (69, 178, 218), (68, 185, 219), (34, 175, 205), (21, 174, 207), (10, 163, 206), (39, 183, 228), (63, 188, 226), (96, 199, 231), (137, 214, 240), (160, 214, 233), (185, 214, 227), (198, 215, 225), (208, 221, 231), (216, 227, 238), (225, 235, 244), (231, 238, 246), (232, 237, 243), (229, 233, 236), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 1), (0, 0, 3), (0, 0, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 3), (200, 210, 220), (197, 210, 225), (197, 211, 227), (197, 212, 226), (200, 212, 224), (201, 214, 225), (199, 214, 227), (198, 215, 226), (197, 214, 222), (203, 218, 224), (203, 214, 222), (209, 214, 216), (218, 215, 201), (231, 213, 173), (250, 211, 132), (255, 203, 86), (252, 184, 30), (255, 181, 17), (255, 169, 20), (255, 160, 28), (255, 144, 32), (253, 129, 33), (238, 108, 24), (204, 69, 7), (177, 39, 9), (157, 17, 3), (154, 12, 0), (200, 54, 39), (218, 62, 46), (220, 61, 47), (215, 60, 51), (184, 40, 14), (181, 56, 0), (196, 80, 0), (222, 106, 29), (224, 108, 51), (161, 44, 26), (144, 32, 36), (129, 26, 39), (126, 29, 46), (131, 34, 51), (142, 38, 56), (165, 44, 69), (182, 51, 77), (188, 50, 75), (173, 47, 70), (156, 61, 82), (105, 46, 69), (31, 15, 45), (15, 23, 62), (24, 36, 87), (22, 48, 105), (11, 60, 116), (6, 71, 129), (7, 79, 143), (18, 95, 164), (35, 117, 191), (55, 144, 218), (43, 145, 212), (25, 134, 193), (52, 165, 214), (99, 205, 245), (137, 227, 255), (117, 212, 241), (79, 198, 222), (46, 183, 210), (17, 165, 201), (20, 172, 211), (18, 166, 203), (31, 162, 197), (51, 154, 187), (110, 183, 208), (183, 221, 234), (219, 238, 246), (225, 238, 247), (224, 234, 243), (228, 237, 245), (227, 235, 241), (227, 234, 238), (234, 238, 242), (0, 0, 3), (1, 0, 1), (1, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (3, 0, 0), (3, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 1), (0, 0, 3), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 3), (200, 210, 220), (196, 211, 225), (196, 211, 227), (197, 211, 227), (201, 212, 224), (200, 212, 223), (198, 214, 226), (198, 215, 226), (201, 217, 225), (201, 215, 223), (202, 212, 222), (208, 213, 218), (217, 216, 210), (237, 224, 189), (255, 226, 144), (255, 210, 83), (255, 200, 29), (251, 184, 1), (254, 178, 14), (252, 163, 20), (232, 126, 7), (234, 115, 19), (226, 97, 21), (171, 37, 0), (155, 20, 0), (156, 20, 12), (149, 12, 0), (174, 28, 11), (195, 33, 22), (196, 26, 25), (191, 24, 34), (201, 46, 42), (205, 73, 26), (225, 106, 41), (216, 100, 42), (184, 70, 33), (155, 42, 37), (133, 27, 42), (106, 12, 34), (117, 28, 51), (130, 40, 59), (141, 40, 61), (168, 48, 74), (178, 47, 73), (189, 54, 77), (203, 81, 102), (182, 90, 110), (101, 46, 70), (40, 28, 60), (6, 18, 59), (6, 22, 74), (8, 38, 93), (3, 57, 110), (0, 69, 123), (0, 74, 135), (5, 86, 152), (9, 93, 162), (16, 109, 177), (22, 127, 190), (21, 132, 189), (42, 153, 202), (68, 172, 215), (101, 192, 230), (117, 207, 241), (109, 214, 242), (67, 184, 211), (34, 159, 190), (15, 147, 179), (23, 162, 192), (13, 141, 171), (9, 107, 142), (91, 159, 188), (154, 192, 206), (204, 223, 230), (225, 237, 246), (226, 234, 244), (226, 235, 242), (227, 235, 241), (228, 236, 240), (227, 232, 236), (0, 0, 4), (1, 0, 3), (0, 0, 1), (0, 0, 0), (0, 1, 0), (0, 0, 0), (4, 0, 0), (4, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 1), (0, 0, 3), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 3), (199, 209, 219), (196, 211, 225), (196, 211, 227), (197, 211, 227), (200, 211, 223), (200, 212, 223), (197, 213, 225), (198, 215, 226), (200, 214, 223), (200, 211, 221), (202, 212, 224), (211, 216, 218), (223, 219, 198), (243, 227, 166), (255, 228, 109), (247, 205, 45), (253, 196, 12), (255, 186, 1), (255, 177, 15), (232, 136, 0), (192, 84, 0), (206, 86, 0), (213, 81, 25), (155, 20, 0), (146, 14, 7), (140, 11, 9), (140, 13, 0), (164, 27, 10), (185, 28, 18), (209, 42, 41), (197, 32, 40), (190, 37, 31), (217, 87, 44), (255, 136, 81), (192, 73, 32), (162, 46, 25), (135, 23, 33), (118, 15, 41), (100, 12, 38), (106, 25, 50), (110, 26, 50), (127, 35, 58), (152, 44, 68), (146, 30, 53), (152, 33, 54), (172, 66, 88), (150, 70, 96), (85, 39, 70), (33, 28, 66), (0, 19, 63), (5, 32, 83), (10, 53, 106), (2, 68, 119), (0, 77, 131), (0, 82, 146), (12, 101, 167), (7, 107, 168), (0, 103, 162), (1, 111, 169), (10, 123, 181), (27, 140, 198), (11, 123, 179), (7, 115, 169), (48, 153, 201), (106, 205, 246), (146, 239, 255), (126, 208, 238), (84, 169, 193), (62, 160, 178), (67, 158, 178), (141, 201, 235), (165, 205, 237), (194, 223, 238), (213, 232, 240), (222, 233, 243), (226, 234, 244), (226, 233, 242), (224, 231, 238), (228, 236, 240), (230, 235, 239), (0, 0, 4), (1, 0, 3), (0, 0, 1), (0, 0, 0), (0, 1, 0), (0, 0, 0), (4, 0, 0), (4, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 1), (0, 0, 3), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 3), (199, 209, 219), (195, 210, 224), (196, 211, 227), (196, 210, 226), (200, 211, 223), (199, 211, 222), (197, 213, 225), (198, 214, 224), (196, 208, 214), (203, 212, 218), (205, 214, 223), (217, 219, 213), (233, 224, 183), (246, 226, 139), (254, 223, 78), (252, 207, 28), (252, 191, 3), (252, 176, 0), (255, 167, 8), (255, 156, 21), (240, 130, 20), (226, 105, 25), (205, 71, 25), (165, 29, 8), (138, 11, 5), (124, 0, 0), (132, 7, 0), (163, 28, 13), (184, 30, 21), (221, 57, 54), (215, 52, 55), (192, 39, 33), (229, 94, 62), (255, 131, 94), (200, 77, 56), (167, 50, 48), (120, 15, 32), (103, 11, 39), (92, 15, 42), (82, 14, 39), (89, 22, 46), (98, 26, 48), (109, 26, 46), (104, 15, 35), (121, 32, 54), (131, 52, 79), (109, 52, 87), (90, 61, 101), (38, 44, 88), (0, 24, 72), (4, 36, 87), (12, 57, 110), (11, 77, 128), (16, 91, 148), (14, 90, 158), (15, 98, 168), (6, 100, 163), (0, 97, 156), (0, 103, 159), (1, 108, 163), (1, 110, 168), (0, 103, 164), (4, 116, 179), (45, 156, 216), (76, 183, 234), (93, 187, 229), (165, 238, 255), (181, 245, 255), (169, 237, 249), (173, 232, 245), (195, 231, 255), (200, 225, 249), (213, 236, 250), (210, 229, 238), (212, 223, 234), (225, 232, 243), (227, 234, 243), (225, 232, 239), (228, 236, 240), (227, 232, 236), (0, 0, 4), (1, 0, 2), (0, 0, 1), (0, 1, 0), (0, 1, 0), (0, 1, 0), (3, 0, 0), (4, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 1), (0, 0, 3), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 4), (199, 209, 220), (195, 209, 225), (195, 210, 226), (196, 210, 226), (199, 210, 222), (199, 211, 223), (196, 212, 225), (197, 213, 222), (202, 212, 213), (209, 216, 215), (207, 213, 214), (219, 218, 198), (240, 224, 159), (243, 214, 102), (242, 204, 41), (249, 198, 12), (249, 180, 0), (255, 172, 1), (255, 156, 2), (242, 134, 0), (235, 123, 13), (232, 111, 30), (206, 71, 24), (164, 28, 4), (136, 15, 1), (127, 7, 0), (123, 0, 0), (166, 25, 15), (203, 47, 39), (215, 53, 47), (209, 50, 46), (221, 67, 60), (212, 66, 51), (209, 71, 60), (216, 85, 91), (158, 43, 59), (113, 21, 41), (90, 17, 38), (73, 12, 35), (64, 15, 37), (56, 16, 35), (55, 15, 32), (62, 15, 30), (58, 8, 26), (68, 19, 45), (73, 33, 68), (62, 39, 85), (76, 72, 123), (44, 63, 114), (3, 33, 84), (4, 34, 85), (5, 42, 94), (6, 57, 111), (24, 81, 142), (20, 77, 149), (12, 72, 149), (14, 80, 156), (6, 82, 150), (3, 90, 146), (2, 96, 148), (0, 90, 144), (4, 102, 160), (18, 120, 187), (5, 116, 182), (14, 142, 199), (41, 163, 210), (108, 204, 239), (170, 240, 255), (198, 245, 255), (199, 230, 240), (204, 228, 237), (206, 227, 236), (202, 224, 232), (206, 225, 234), (214, 225, 236), (219, 226, 237), (216, 223, 232), (220, 227, 234), (228, 236, 240), (225, 230, 234), (0, 0, 3), (1, 0, 2), (0, 0, 1), (0, 1, 0), (0, 2, 0), (0, 1, 0), (2, 0, 0), (3, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 1), (0, 0, 3), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 4), (198, 208, 219), (195, 209, 225), (195, 209, 226), (195, 209, 225), (199, 210, 223), (198, 210, 222), (195, 211, 224), (197, 212, 223), (203, 212, 215), (211, 216, 212), (210, 212, 203), (228, 220, 181), (249, 226, 132), (243, 207, 69), (237, 189, 18), (241, 179, 0), (253, 175, 5), (248, 155, 0), (255, 150, 4), (251, 138, 8), (232, 117, 9), (223, 101, 18), (209, 74, 17), (181, 47, 10), (139, 20, 0), (128, 9, 0), (145, 10, 0), (203, 56, 47), (228, 71, 63), (201, 41, 32), (199, 41, 30), (239, 84, 73), (231, 80, 71), (223, 80, 81), (221, 92, 112), (161, 52, 80), (114, 33, 58), (76, 17, 40), (51, 7, 30), (46, 14, 35), (41, 17, 34), (40, 17, 33), (50, 23, 39), (39, 13, 35), (24, 4, 39), (32, 22, 69), (33, 38, 95), (45, 64, 124), (37, 69, 124), (3, 40, 91), (8, 41, 90), (2, 38, 87), (1, 46, 100), (26, 76, 136), (20, 71, 140), (5, 57, 130), (14, 68, 141), (21, 83, 150), (9, 85, 140), (8, 91, 141), (0, 84, 136), (0, 84, 142), (8, 101, 169), (11, 118, 187), (13, 143, 203), (19, 152, 201), (47, 161, 198), (101, 191, 217), (164, 224, 240), (205, 243, 252), (210, 235, 240), (215, 234, 239), (213, 234, 242), (214, 232, 242), (217, 228, 239), (221, 228, 239), (214, 221, 230), (213, 220, 227), (225, 233, 237), (230, 235, 238), (0, 0, 3), (1, 0, 1), (0, 0, 0), (0, 1, 0), (0, 2, 0), (0, 1, 0), (2, 0, 0), (3, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 2), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 4), (198, 208, 219), (194, 208, 224), (194, 208, 226), (195, 209, 226), (198, 209, 223), (198, 210, 223), (195, 211, 225), (196, 211, 224), (199, 207, 218), (206, 208, 207), (219, 214, 193), (240, 225, 161), (252, 221, 95), (250, 205, 43), (252, 192, 20), (250, 176, 7), (247, 159, 7), (245, 145, 4), (255, 147, 11), (244, 129, 5), (226, 109, 5), (237, 113, 24), (233, 102, 22), (203, 73, 14), (138, 18, 0), (125, 1, 0), (175, 33, 19), (217, 64, 50), (203, 47, 35), (180, 22, 10), (205, 46, 29), (242, 85, 67), (222, 70, 55), (221, 82, 79), (178, 57, 79), (144, 46, 80), (105, 32, 68), (64, 14, 48), (41, 14, 41), (32, 14, 36), (33, 13, 32), (29, 7, 28), (30, 7, 32), (23, 7, 42), (13, 9, 60), (24, 35, 98), (23, 50, 120), (28, 67, 134), (31, 76, 132), (0, 45, 93), (10, 51, 95), (5, 47, 90), (6, 55, 103), (33, 87, 140), (18, 77, 134), (0, 52, 110), (0, 58, 114), (4, 65, 119), (0, 70, 120), (7, 84, 135), (10, 89, 144), (5, 88, 147), (0, 83, 148), (0, 93, 158), (4, 120, 179), (20, 144, 195), (31, 157, 196), (45, 165, 191), (86, 192, 207), (155, 232, 242), (200, 236, 250), (210, 228, 241), (214, 235, 246), (210, 228, 239), (215, 226, 238), (227, 234, 246), (226, 233, 242), (218, 225, 232), (223, 231, 235), (228, 233, 236), (0, 0, 3), (1, 0, 1), (0, 0, 0), (0, 1, 0), (0, 2, 0), (0, 2, 0), (1, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 2), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 4), (198, 208, 219), (194, 208, 225), (194, 208, 226), (195, 209, 226), (198, 209, 223), (197, 209, 222), (195, 211, 225), (196, 211, 225), (205, 213, 228), (208, 208, 208), (226, 216, 183), (239, 218, 137), (233, 196, 55), (237, 185, 14), (253, 184, 14), (250, 166, 7), (245, 150, 8), (247, 143, 11), (255, 149, 18), (246, 132, 11), (220, 101, 1), (216, 93, 4), (219, 92, 4), (217, 91, 22), (157, 38, 4), (128, 4, 0), (166, 26, 10), (169, 20, 7), (152, 4, 0), (174, 24, 11), (219, 65, 45), (238, 87, 66), (196, 56, 41), (184, 59, 59), (144, 40, 65), (115, 30, 69), (103, 35, 77), (60, 15, 54), (32, 17, 47), (13, 9, 34), (19, 7, 29), (25, 10, 34), (22, 8, 40), (21, 17, 60), (18, 29, 88), (18, 44, 113), (21, 62, 135), (50, 100, 168), (22, 73, 128), (2, 53, 99), (21, 68, 110), (10, 58, 100), (0, 49, 95), (17, 74, 124), (11, 71, 121), (0, 55, 103), (1, 60, 104), (0, 55, 99), (7, 78, 125), (9, 85, 136), (0, 71, 126), (22, 106, 163), (18, 111, 168), (0, 85, 140), (0, 79, 132), (17, 130, 178), (28, 149, 189), (37, 162, 194), (50, 173, 195), (84, 185, 204), (161, 220, 243), (202, 236, 255), (207, 233, 248), (216, 235, 247), (220, 232, 245), (224, 232, 244), (225, 232, 242), (225, 232, 239), (228, 236, 240), (226, 231, 234), (0, 0, 3), (1, 0, 1), (0, 0, 0), (0, 1, 0), (0, 2, 0), (0, 2, 0), (1, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 2), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 4), (198, 208, 219), (194, 208, 225), (194, 208, 226), (194, 208, 225), (197, 208, 222), (196, 208, 221), (194, 210, 225), (195, 209, 226), (201, 210, 227), (206, 205, 203), (226, 212, 168), (232, 204, 115), (222, 180, 42), (241, 184, 20), (245, 170, 7), (243, 154, 0), (240, 141, 3), (238, 134, 3), (247, 142, 10), (255, 146, 26), (203, 86, 0), (195, 73, 0), (218, 96, 14), (206, 86, 17), (169, 53, 10), (139, 20, 0), (156, 25, 11), (152, 16, 9), (132, 0, 0), (179, 44, 34), (234, 91, 72), (203, 66, 48), (149, 31, 25), (108, 9, 19), (97, 19, 49), (108, 41, 82), (107, 40, 83), (61, 15, 54), (19, 12, 45), (8, 16, 44), (6, 6, 30), (17, 14, 41), (12, 12, 47), (21, 31, 76), (31, 54, 114), (25, 60, 127), (30, 76, 143), (48, 99, 161), (24, 73, 124), (2, 52, 97), (12, 64, 107), (14, 68, 113), (2, 58, 108), (0, 53, 104), (4, 59, 107), (0, 56, 99), (3, 63, 99), (0, 64, 101), (16, 89, 133), (22, 101, 151), (37, 120, 173), (37, 127, 179), (21, 124, 167), (6, 112, 152), (0, 95, 135), (0, 86, 128), (0, 98, 142), (15, 118, 161), (17, 131, 168), (47, 157, 191), (58, 151, 185), (136, 206, 234), (206, 245, 255), (211, 231, 242), (220, 232, 245), (219, 227, 239), (219, 226, 236), (227, 234, 242), (226, 234, 239), (225, 230, 233), (0, 0, 3), (1, 0, 1), (0, 0, 0), (0, 1, 0), (0, 2, 0), (0, 2, 0), (1, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 2), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 4), (197, 207, 218), (193, 207, 224), (193, 207, 225), (193, 207, 225), (196, 207, 221), (196, 208, 222), (193, 209, 224), (195, 210, 226), (199, 209, 225), (204, 205, 198), (227, 212, 161), (231, 202, 111), (232, 190, 65), (242, 184, 39), (242, 167, 14), (230, 142, 0), (218, 120, 0), (230, 128, 2), (239, 138, 12), (245, 141, 27), (210, 97, 9), (188, 73, 0), (191, 80, 7), (181, 73, 10), (161, 57, 11), (153, 47, 16), (151, 35, 20), (149, 31, 26), (120, 7, 8), (177, 61, 62), (186, 61, 54), (138, 20, 15), (109, 15, 22), (76, 4, 23), (75, 22, 56), (107, 59, 101), (101, 42, 88), (72, 28, 71), (14, 13, 45), (1, 17, 43), (14, 24, 50), (0, 8, 38), (1, 11, 49), (1, 18, 64), (5, 34, 90), (21, 60, 119), (5, 51, 108), (2, 50, 103), (24, 69, 116), (11, 61, 105), (20, 81, 126), (13, 79, 128), (3, 70, 123), (11, 75, 127), (8, 65, 112), (0, 45, 87), (0, 50, 89), (12, 78, 118), (16, 90, 134), (5, 84, 131), (106, 187, 234), (97, 183, 226), (40, 136, 169), (1, 98, 127), (30, 119, 151), (48, 133, 169), (63, 149, 191), (19, 112, 156), (0, 99, 142), (0, 90, 131), (16, 123, 161), (70, 156, 187), (166, 211, 230), (215, 236, 248), (217, 229, 243), (223, 231, 244), (229, 236, 247), (228, 235, 243), (220, 228, 233), (225, 230, 233), (0, 0, 3), (1, 0, 1), (0, 0, 0), (0, 1, 0), (0, 2, 0), (0, 2, 0), (1, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 2), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 4), (196, 206, 217), (192, 206, 223), (192, 206, 224), (192, 206, 224), (196, 207, 222), (195, 207, 221), (193, 209, 224), (193, 209, 223), (203, 216, 226), (205, 209, 195), (224, 213, 157), (244, 218, 134), (254, 216, 118), (254, 201, 84), (237, 169, 28), (219, 138, 0), (215, 123, 0), (203, 106, 0), (215, 120, 4), (221, 122, 19), (182, 78, 0), (175, 71, 6), (208, 112, 53), (205, 117, 64), (141, 60, 15), (137, 53, 19), (206, 111, 92), (174, 78, 73), (117, 27, 38), (126, 35, 52), (131, 30, 47), (118, 25, 43), (98, 30, 52), (60, 13, 41), (50, 21, 58), (68, 39, 84), (102, 55, 108), (66, 29, 75), (5, 7, 33), (3, 23, 43), (4, 20, 48), (0, 13, 49), (9, 24, 65), (1, 21, 66), (0, 16, 64), (9, 44, 91), (5, 45, 88), (0, 29, 70), (0, 40, 82), (18, 69, 113), (29, 103, 150), (6, 90, 141), (0, 75, 129), (0, 77, 130), (0, 65, 112), (0, 53, 100), (0, 57, 109), (8, 74, 126), (11, 86, 132), (48, 125, 166), (113, 186, 221), (116, 187, 217), (122, 194, 218), (94, 166, 189), (105, 176, 203), (108, 184, 215), (101, 188, 222), (80, 174, 211), (31, 126, 166), (43, 141, 181), (45, 146, 184), (52, 135, 166), (131, 175, 194), (200, 221, 234), (203, 216, 230), (218, 227, 240), (217, 225, 236), (223, 230, 238), (228, 236, 241), (226, 231, 234), (0, 0, 3), (1, 0, 1), (0, 0, 0), (0, 1, 0), (0, 2, 0), (0, 1, 0), (1, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 2), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 5), (195, 205, 217), (191, 205, 222), (191, 205, 224), (191, 205, 223), (195, 205, 221), (195, 207, 222), (193, 209, 225), (194, 210, 224), (196, 210, 219), (202, 209, 196), (203, 197, 146), (224, 206, 134), (239, 209, 133), (255, 218, 125), (242, 185, 64), (227, 156, 29), (207, 123, 8), (197, 106, 0), (192, 100, 0), (194, 100, 11), (168, 74, 2), (174, 85, 26), (216, 141, 90), (249, 185, 141), (192, 134, 96), (178, 117, 90), (201, 126, 114), (154, 75, 78), (97, 24, 43), (114, 40, 67), (101, 21, 48), (105, 33, 61), (95, 44, 75), (53, 22, 56), (46, 33, 69), (45, 32, 75), (96, 66, 119), (63, 40, 87), (11, 20, 44), (2, 26, 45), (1, 26, 55), (10, 34, 71), (5, 26, 70), (4, 28, 73), (0, 28, 71), (2, 42, 82), (21, 66, 99), (0, 29, 62), (1, 43, 82), (23, 77, 120), (50, 131, 177), (9, 102, 151), (5, 97, 148), (43, 126, 176), (42, 112, 156), (12, 76, 122), (9, 74, 131), (5, 75, 130), (83, 163, 206), (142, 220, 255), (134, 198, 226), (157, 212, 235), (156, 207, 226), (165, 215, 234), (160, 211, 233), (148, 205, 230), (117, 185, 213), (84, 159, 189), (83, 160, 194), (93, 176, 211), (76, 167, 201), (107, 185, 213), (173, 217, 235), (210, 232, 246), (196, 211, 225), (217, 226, 240), (224, 232, 243), (219, 228, 235), (223, 231, 236), (225, 230, 233), (0, 0, 3), (1, 0, 1), (0, 0, 0), (0, 1, 0), (0, 2, 0), (0, 1, 0), (1, 0, 0), (2, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 2), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 5), (194, 204, 216), (190, 204, 222), (191, 205, 225), (191, 205, 224), (195, 205, 222), (195, 207, 222), (193, 209, 225), (194, 210, 225), (194, 208, 220), (208, 217, 213), (197, 200, 164), (195, 189, 135), (203, 187, 129), (231, 203, 132), (222, 180, 87), (208, 150, 49), (211, 136, 38), (199, 113, 22), (176, 84, 2), (166, 76, 3), (132, 51, 0), (157, 89, 34), (196, 147, 99), (228, 190, 152), (192, 162, 137), (209, 171, 161), (165, 107, 114), (115, 48, 67), (98, 34, 60), (90, 27, 55), (96, 32, 56), (118, 61, 86), (91, 51, 84), (47, 24, 59), (47, 43, 76), (32, 33, 70), (34, 27, 73), (27, 26, 69), (7, 25, 52), (0, 14, 36), (0, 37, 65), (17, 54, 90), (0, 30, 75), (0, 31, 79), (4, 46, 89), (0, 47, 84), (25, 84, 114), (0, 52, 83), (0, 37, 75), (17, 77, 119), (24, 107, 149), (5, 98, 141), (27, 117, 160), (87, 169, 211), (117, 189, 229), (12, 79, 123), (4, 74, 128), (5, 82, 135), (50, 140, 177), (102, 184, 213), (157, 210, 236), (177, 215, 237), (165, 200, 217), (194, 226, 241), (194, 222, 240), (190, 217, 236), (179, 208, 230), (148, 184, 207), (149, 199, 223), (106, 169, 194), (65, 144, 168), (77, 148, 169), (121, 163, 178), (184, 207, 221), (191, 206, 220), (196, 207, 220), (221, 231, 241), (223, 232, 239), (220, 228, 233), (229, 234, 237), (0, 0, 3), (2, 0, 1), (1, 0, 0), (0, 1, 0), (0, 2, 0), (0, 1, 0), (1, 0, 1), (2, 0, 1), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 2), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 5), (194, 203, 217), (190, 204, 222), (191, 205, 225), (191, 205, 224), (195, 205, 222), (195, 207, 222), (193, 209, 225), (194, 210, 226), (193, 206, 221), (202, 213, 216), (204, 214, 195), (200, 205, 172), (213, 209, 171), (217, 202, 155), (231, 201, 142), (234, 187, 115), (179, 114, 25), (172, 93, 1), (169, 80, 0), (174, 89, 17), (142, 72, 10), (192, 142, 91), (221, 192, 153), (212, 196, 172), (201, 190, 180), (196, 175, 180), (121, 78, 97), (90, 33, 60), (88, 26, 58), (103, 40, 71), (104, 43, 68), (112, 61, 86), (85, 48, 81), (41, 22, 56), (49, 49, 78), (26, 35, 67), (8, 18, 59), (7, 25, 63), (30, 62, 84), (28, 72, 89), (0, 47, 70), (14, 66, 98), (6, 46, 92), (0, 39, 90), (4, 58, 104), (0, 64, 103), (26, 107, 137), (29, 108, 138), (0, 51, 90), (0, 54, 95), (24, 105, 143), (22, 107, 143), (84, 163, 197), (146, 219, 253), (106, 175, 209), (9, 78, 117), (16, 92, 140), (30, 111, 157), (19, 105, 138), (61, 134, 160), (159, 199, 224), (209, 233, 253), (207, 232, 245), (211, 232, 243), (216, 230, 241), (215, 225, 237), (207, 218, 231), (217, 236, 249), (194, 227, 241), (159, 206, 222), (125, 185, 202), (95, 152, 169), (117, 155, 169), (184, 209, 222), (213, 229, 243), (206, 217, 230), (214, 224, 234), (222, 231, 238), (222, 230, 235), (224, 229, 232), (1, 0, 3), (2, 0, 1), (1, 0, 0), (0, 0, 0), (0, 1, 0), (0, 1, 0), (1, 0, 1), (2, 0, 1), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 2), (0, 1, 2), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 5), (194, 203, 217), (190, 204, 222), (190, 204, 224), (191, 205, 224), (195, 205, 222), (195, 207, 222), (193, 209, 226), (193, 209, 226), (200, 212, 227), (193, 205, 216), (194, 210, 211), (192, 206, 199), (203, 210, 193), (194, 189, 169), (219, 199, 181), (238, 202, 161), (222, 168, 80), (219, 148, 41), (197, 112, 13), (179, 99, 13), (156, 98, 31), (200, 165, 119), (208, 194, 173), (195, 194, 190), (198, 198, 205), (173, 163, 180), (160, 129, 153), (128, 79, 109), (149, 83, 119), (182, 109, 145), (183, 113, 145), (143, 84, 115), (98, 59, 92), (80, 61, 92), (96, 95, 120), (63, 77, 104), (17, 39, 77), (0, 33, 65), (33, 83, 93), (52, 114, 117), (18, 89, 101), (25, 92, 118), (6, 57, 103), (2, 53, 108), (3, 73, 125), (5, 93, 139), (21, 128, 163), (36, 140, 174), (7, 87, 128), (0, 54, 95), (24, 96, 129), (78, 147, 175), (147, 207, 232), (171, 230, 254), (103, 164, 191), (28, 97, 129), (0, 80, 118), (27, 108, 146), (36, 105, 137), (149, 199, 227), (195, 219, 245), (199, 214, 233), (215, 235, 244), (210, 228, 232), (220, 227, 231), (229, 234, 238), (216, 229, 231), (213, 233, 235), (211, 239, 243), (189, 222, 229), (183, 220, 230), (160, 196, 209), (193, 225, 238), (200, 225, 239), (207, 225, 238), (220, 232, 245), (216, 227, 237), (218, 227, 234), (223, 231, 236), (226, 231, 234), (1, 0, 3), (2, 0, 1), (1, 0, 0), (0, 0, 0), (0, 1, 0), (0, 1, 0), (2, 0, 1), (3, 0, 1), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 2), (0, 0, 2), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 1, 5), (194, 203, 217), (191, 204, 223), (189, 204, 223), (191, 205, 223), (193, 206, 222), (194, 207, 223), (194, 208, 226), (194, 208, 225), (197, 207, 221), (199, 210, 223), (195, 213, 226), (195, 213, 223), (201, 215, 217), (200, 205, 206), (217, 209, 214), (223, 201, 184), (201, 164, 96), (177, 126, 36), (167, 103, 18), (158, 98, 25), (135, 97, 42), (185, 166, 133), (210, 210, 202), (190, 200, 208), (188, 200, 215), (179, 183, 203), (180, 165, 188), (184, 148, 176), (167, 110, 144), (196, 129, 164), (207, 139, 172), (193, 134, 165), (122, 80, 111), (144, 120, 146), (165, 159, 177), (130, 139, 154), (20, 43, 62), (19, 56, 66), (58, 108, 97), (74, 136, 121), (59, 132, 132), (57, 128, 148), (14, 74, 117), (8, 72, 126), (0, 79, 132), (0, 99, 146), (9, 128, 166), (23, 140, 175), (32, 124, 164), (0, 68, 105), (28, 96, 124), (118, 177, 198), (146, 193, 209), (174, 217, 234), (181, 227, 251), (137, 191, 219), (52, 119, 148), (97, 163, 192), (154, 204, 231), (184, 217, 242), (178, 194, 217), (211, 222, 239), (206, 223, 230), (218, 233, 236), (224, 229, 232), (221, 225, 227), (224, 236, 235), (215, 232, 232), (211, 232, 234), (210, 232, 236), (216, 236, 244), (195, 216, 226), (197, 220, 230), (213, 234, 245), (208, 223, 235), (222, 233, 244), (218, 229, 238), (224, 233, 240), (223, 231, 236), (227, 232, 235), (0, 0, 3), (1, 0, 1), (1, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (2, 0, 1), (2, 0, 1), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 2), (1, 0, 2), (2, 0, 1), (1, 0, 0), (0, 1, 0), (0, 1, 4), (193, 202, 218), (190, 202, 223), (187, 204, 221), (188, 206, 221), (190, 206, 222), (192, 207, 223), (193, 207, 225), (196, 208, 223), (201, 208, 219), (200, 208, 219), (196, 209, 225), (193, 210, 228), (194, 211, 229), (196, 211, 226), (203, 210, 222), (210, 209, 207), (217, 206, 179), (178, 159, 119), (152, 126, 85), (126, 102, 66), (132, 119, 94), (199, 197, 185), (211, 219, 223), (189, 206, 218), (171, 195, 208), (188, 207, 222), (187, 190, 208), (207, 191, 212), (194, 159, 184), (158, 109, 137), (159, 104, 133), (146, 93, 121), (144, 100, 125), (191, 159, 178), (186, 169, 176), (152, 150, 146), (115, 126, 113), (104, 127, 100), (79, 112, 69), (110, 155, 116), (78, 135, 123), (70, 135, 147), (22, 90, 125), (15, 93, 139), (2, 97, 144), (0, 96, 140), (9, 127, 164), (22, 138, 172), (41, 141, 178), (45, 130, 163), (99, 169, 191), (117, 172, 185), (137, 176, 184), (187, 215, 227), (198, 218, 243), (202, 223, 252), (192, 224, 246), (198, 233, 252), (199, 228, 245), (189, 212, 228), (179, 195, 210), (204, 216, 229), (218, 232, 240), (217, 230, 236), (221, 229, 234), (222, 229, 235), (223, 232, 237), (221, 232, 237), (219, 231, 236), (218, 230, 236), (218, 230, 237), (219, 230, 238), (213, 225, 232), (212, 222, 229), (217, 226, 233), (222, 231, 238), (222, 231, 238), (221, 230, 236), (224, 230, 235), (226, 231, 234), (0, 0, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (193, 202, 219), (190, 202, 224), (187, 204, 220), (187, 206, 220), (189, 207, 222), (191, 207, 223), (193, 207, 224), (197, 208, 223), (201, 208, 218), (201, 208, 219), (196, 209, 225), (193, 210, 230), (191, 211, 234), (192, 211, 232), (197, 212, 226), (202, 211, 217), (211, 213, 209), (216, 214, 202), (220, 215, 201), (199, 195, 182), (195, 196, 189), (211, 218, 219), (185, 198, 208), (159, 178, 192), (167, 192, 205), (175, 196, 209), (186, 195, 210), (212, 207, 226), (223, 204, 225), (148, 117, 141), (111, 74, 100), (131, 93, 118), (190, 156, 178), (181, 155, 169), (196, 181, 184), (160, 156, 145), (91, 97, 70), (88, 102, 60), (83, 103, 48), (116, 145, 96), (82, 123, 97), (94, 147, 145), (33, 96, 117), (14, 90, 124), (0, 89, 127), (0, 98, 137), (18, 128, 163), (16, 124, 159), (44, 142, 180), (88, 172, 207), (125, 194, 216), (137, 189, 202), (140, 176, 181), (190, 213, 221), (200, 212, 235), (210, 219, 245), (201, 217, 234), (202, 220, 233), (207, 225, 237), (209, 226, 237), (200, 215, 226), (206, 220, 230), (213, 226, 234), (213, 225, 232), (217, 227, 234), (220, 229, 236), (223, 230, 238), (223, 230, 237), (222, 229, 236), (221, 228, 235), (221, 228, 235), (223, 229, 236), (223, 229, 234), (220, 226, 231), (223, 229, 235), (226, 234, 240), (223, 232, 238), (223, 231, 237), (225, 231, 236), (226, 231, 234), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (193, 202, 219), (190, 202, 224), (187, 204, 220), (187, 206, 220), (189, 207, 222), (191, 207, 223), (193, 207, 224), (196, 208, 223), (199, 209, 220), (198, 209, 220), (195, 210, 224), (193, 212, 228), (192, 212, 229), (193, 213, 229), (197, 212, 224), (201, 213, 219), (209, 215, 215), (208, 209, 205), (217, 215, 211), (218, 217, 214), (211, 215, 216), (171, 180, 185), (140, 154, 165), (166, 182, 196), (192, 207, 220), (153, 164, 178), (197, 200, 216), (216, 213, 231), (204, 194, 214), (146, 131, 153), (131, 114, 138), (154, 139, 162), (161, 150, 171), (180, 175, 189), (191, 192, 196), (179, 184, 176), (99, 107, 85), (136, 146, 111), (119, 129, 83), (111, 126, 78), (161, 186, 146), (119, 154, 130), (87, 132, 134), (84, 142, 160), (58, 132, 158), (34, 120, 151), (32, 126, 159), (44, 138, 175), (49, 136, 179), (73, 150, 191), (123, 188, 217), (153, 206, 223), (155, 195, 202), (192, 222, 229), (194, 214, 231), (208, 225, 245), (206, 222, 237), (202, 219, 231), (208, 225, 236), (214, 229, 240), (212, 226, 236), (210, 223, 232), (215, 226, 235), (215, 225, 233), (216, 225, 232), (218, 227, 234), (222, 230, 236), (223, 230, 237), (223, 230, 237), (222, 229, 236), (222, 229, 236), (223, 229, 235), (225, 231, 236), (222, 228, 233), (223, 229, 235), (225, 233, 239), (222, 231, 237), (222, 230, 236), (224, 230, 235), (225, 230, 233), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (193, 202, 219), (190, 202, 224), (187, 204, 220), (187, 206, 220), (189, 207, 222), (191, 207, 223), (193, 207, 224), (194, 207, 223), (197, 209, 222), (196, 210, 221), (195, 212, 224), (193, 212, 225), (192, 213, 225), (194, 214, 225), (196, 213, 223), (200, 213, 221), (207, 215, 220), (205, 210, 215), (208, 210, 215), (205, 208, 215), (211, 218, 226), (177, 188, 198), (160, 175, 187), (198, 214, 228), (207, 219, 232), (201, 209, 223), (208, 211, 227), (221, 221, 238), (213, 211, 230), (170, 168, 188), (192, 191, 213), (192, 193, 215), (192, 197, 217), (186, 195, 210), (196, 208, 214), (154, 166, 162), (105, 116, 100), (169, 178, 151), (150, 156, 120), (142, 152, 110), (156, 174, 132), (135, 162, 131), (159, 194, 187), (143, 189, 197), (122, 181, 198), (119, 188, 212), (101, 176, 204), (90, 166, 199), (112, 181, 223), (106, 168, 209), (119, 173, 203), (163, 208, 228), (195, 234, 241), (189, 221, 226), (200, 225, 238), (198, 218, 234), (210, 226, 240), (209, 224, 236), (213, 228, 239), (209, 223, 233), (212, 225, 234), (214, 225, 235), (222, 232, 241), (219, 229, 237), (217, 226, 233), (220, 228, 234), (222, 230, 235), (223, 230, 236), (222, 229, 235), (222, 229, 235), (222, 229, 235), (223, 229, 235), (224, 230, 235), (221, 227, 232), (222, 228, 234), (223, 231, 237), (220, 229, 235), (221, 229, 235), (224, 230, 235), (224, 229, 232), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (192, 201, 218), (190, 202, 224), (187, 204, 220), (187, 206, 220), (189, 207, 222), (191, 207, 223), (193, 207, 224), (193, 207, 224), (195, 210, 224), (194, 211, 223), (193, 211, 221), (194, 213, 222), (193, 213, 221), (195, 214, 222), (196, 213, 222), (199, 213, 223), (200, 211, 222), (204, 213, 226), (209, 215, 230), (201, 208, 224), (210, 220, 235), (199, 212, 226), (189, 205, 218), (202, 219, 231), (202, 216, 229), (211, 222, 235), (209, 218, 233), (205, 211, 227), (210, 216, 233), (201, 207, 225), (199, 207, 227), (196, 207, 227), (199, 214, 233), (200, 217, 233), (189, 207, 217), (159, 177, 179), (116, 132, 123), (173, 186, 168), (168, 178, 152), (152, 164, 134), (149, 170, 139), (159, 187, 164), (166, 198, 194), (161, 198, 206), (141, 186, 199), (138, 188, 205), (144, 196, 217), (147, 197, 223), (154, 198, 233), (146, 186, 221), (136, 171, 198), (137, 169, 186), (201, 231, 237), (206, 234, 237), (198, 224, 233), (210, 232, 245), (207, 223, 236), (212, 226, 237), (218, 232, 242), (212, 225, 234), (216, 227, 237), (218, 228, 237), (223, 233, 241), (218, 227, 234), (220, 228, 234), (221, 229, 234), (221, 229, 234), (222, 229, 235), (221, 228, 234), (222, 229, 235), (222, 229, 235), (224, 230, 236), (224, 230, 235), (222, 228, 233), (223, 229, 235), (223, 231, 237), (221, 230, 236), (222, 230, 236), (225, 231, 236), (225, 230, 233), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (192, 201, 218), (190, 202, 224), (187, 204, 220), (187, 206, 220), (189, 207, 222), (191, 207, 223), (193, 207, 224), (193, 207, 224), (192, 210, 224), (192, 210, 222), (193, 211, 221), (195, 213, 220), (195, 213, 219), (196, 213, 220), (197, 213, 221), (197, 212, 224), (204, 217, 233), (197, 210, 228), (202, 213, 234), (201, 213, 234), (204, 217, 236), (200, 215, 231), (198, 215, 228), (204, 222, 234), (203, 219, 233), (201, 217, 231), (201, 214, 229), (210, 222, 236), (198, 208, 223), (200, 211, 226), (211, 224, 240), (197, 213, 229), (201, 220, 236), (200, 220, 235), (193, 215, 226), (200, 222, 227), (196, 216, 214), (135, 153, 145), (154, 169, 156), (154, 171, 155), (165, 190, 175), (141, 170, 161), (167, 198, 202), (179, 211, 223), (145, 180, 192), (185, 221, 234), (184, 219, 233), (166, 197, 216), (180, 206, 233), (202, 223, 252), (178, 197, 220), (171, 190, 205), (205, 225, 231), (206, 227, 231), (210, 231, 241), (206, 225, 238), (211, 225, 236), (214, 225, 236), (218, 229, 239), (218, 229, 239), (220, 230, 239), (218, 227, 235), (219, 228, 235), (221, 229, 235), (222, 230, 235), (222, 229, 235), (221, 229, 234), (221, 229, 234), (221, 228, 234), (221, 229, 234), (222, 230, 235), (222, 230, 235), (224, 230, 235), (222, 228, 233), (223, 229, 235), (223, 231, 237), (220, 229, 235), (221, 229, 235), (224, 230, 235), (223, 228, 231), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (192, 201, 218), (189, 201, 223), (187, 204, 220), (187, 206, 220), (188, 206, 221), (191, 207, 223), (193, 207, 224), (193, 208, 224), (190, 209, 223), (191, 211, 222), (193, 211, 221), (195, 211, 219), (197, 212, 218), (198, 213, 219), (198, 212, 222), (197, 212, 225), (196, 211, 230), (195, 210, 232), (199, 214, 237), (198, 214, 236), (195, 211, 230), (203, 219, 235), (204, 221, 233), (199, 217, 229), (200, 221, 236), (193, 214, 230), (207, 226, 240), (205, 221, 234), (198, 212, 224), (203, 214, 226), (194, 205, 216), (205, 219, 230), (202, 218, 231), (204, 222, 234), (202, 223, 234), (188, 211, 219), (186, 209, 214), (178, 201, 203), (172, 194, 193), (198, 222, 223), (185, 215, 221), (172, 204, 216), (150, 181, 200), (176, 207, 226), (182, 212, 226), (195, 223, 233), (202, 226, 234), (196, 214, 225), (193, 204, 223), (205, 213, 234), (216, 222, 239), (216, 222, 236), (212, 221, 228), (215, 226, 234), (213, 225, 238), (210, 223, 237), (217, 228, 239), (217, 228, 237), (216, 226, 235), (220, 229, 238), (219, 227, 236), (220, 227, 235), (218, 226, 232), (223, 231, 236), (221, 229, 234), (221, 229, 234), (221, 229, 233), (221, 229, 233), (221, 229, 234), (221, 229, 234), (221, 229, 234), (221, 229, 234), (223, 229, 234), (221, 227, 232), (223, 229, 235), (222, 230, 236), (219, 228, 234), (220, 228, 234), (222, 228, 233), (221, 226, 229), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (192, 201, 218), (189, 201, 223), (187, 204, 220), (186, 205, 219), (188, 206, 221), (191, 207, 223), (192, 206, 223), (193, 208, 224), (190, 209, 223), (190, 210, 221), (193, 210, 220), (196, 210, 220), (198, 211, 219), (199, 211, 220), (199, 211, 223), (198, 211, 226), (199, 214, 233), (195, 212, 233), (195, 213, 234), (200, 218, 238), (194, 211, 229), (201, 218, 233), (203, 218, 230), (202, 219, 231), (197, 217, 233), (197, 218, 235), (199, 218, 233), (201, 218, 230), (203, 217, 227), (205, 218, 226), (206, 218, 225), (208, 221, 229), (206, 222, 230), (203, 221, 231), (211, 231, 241), (182, 203, 214), (164, 186, 197), (213, 236, 245), (203, 225, 235), (199, 223, 235), (191, 218, 235), (147, 175, 196), (187, 215, 238), (183, 210, 231), (176, 201, 215), (199, 222, 231), (202, 221, 226), (213, 226, 233), (199, 207, 220), (214, 217, 234), (219, 221, 236), (223, 224, 237), (220, 223, 232), (214, 219, 229), (218, 224, 238), (218, 226, 240), (218, 227, 237), (222, 231, 239), (217, 226, 234), (220, 227, 236), (218, 225, 233), (223, 230, 237), (220, 226, 232), (221, 227, 233), (220, 226, 232), (221, 227, 232), (220, 228, 232), (221, 229, 233), (222, 230, 235), (222, 230, 235), (220, 229, 234), (220, 228, 233), (222, 228, 233), (221, 227, 232), (223, 229, 235), (222, 230, 236), (220, 229, 235), (221, 229, 235), (223, 229, 234), (222, 227, 230), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (190, 199, 216), (189, 201, 223), (187, 204, 220), (187, 206, 220), (189, 207, 222), (190, 206, 222), (191, 205, 222), (192, 207, 223), (191, 209, 222), (191, 209, 221), (194, 209, 221), (197, 209, 222), (199, 208, 221), (200, 209, 223), (199, 209, 224), (199, 211, 227), (198, 212, 230), (196, 213, 231), (196, 215, 231), (196, 215, 230), (198, 216, 229), (200, 217, 228), (203, 217, 228), (203, 217, 229), (198, 214, 230), (201, 217, 234), (206, 222, 237), (201, 216, 228), (196, 209, 218), (206, 219, 226), (213, 227, 232), (204, 219, 224), (204, 221, 228), (204, 223, 231), (206, 224, 235), (193, 212, 224), (195, 213, 227), (206, 223, 239), (198, 214, 231), (189, 205, 223), (198, 215, 233), (174, 191, 210), (187, 205, 226), (189, 209, 227), (199, 220, 232), (199, 220, 229), (208, 228, 234), (208, 225, 233), (213, 225, 238), (215, 224, 240), (217, 223, 239), (219, 224, 238), (220, 224, 235), (221, 224, 235), (220, 222, 236), (219, 223, 236), (219, 226, 235), (219, 226, 234), (220, 227, 235), (220, 227, 235), (220, 227, 234), (222, 228, 234), (222, 228, 233), (222, 228, 233), (221, 227, 232), (221, 227, 232), (221, 228, 231), (220, 228, 232), (220, 228, 233), (220, 228, 233), (219, 228, 233), (220, 228, 233), (221, 227, 232), (222, 228, 233), (222, 228, 234), (221, 229, 235), (220, 229, 235), (221, 229, 235), (222, 228, 233), (223, 228, 231), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (191, 200, 217), (189, 201, 223), (187, 204, 220), (187, 206, 220), (188, 206, 221), (190, 206, 222), (192, 206, 223), (192, 206, 222), (192, 208, 221), (193, 208, 221), (195, 207, 221), (197, 207, 223), (199, 208, 224), (200, 207, 224), (200, 209, 226), (199, 209, 226), (199, 212, 228), (197, 213, 227), (197, 215, 227), (197, 215, 226), (198, 216, 226), (201, 217, 226), (203, 217, 227), (204, 216, 228), (206, 218, 233), (205, 217, 232), (205, 217, 231), (198, 211, 222), (192, 205, 214), (203, 216, 224), (212, 226, 233), (208, 223, 229), (210, 226, 233), (206, 223, 232), (201, 218, 229), (188, 204, 218), (190, 205, 220), (203, 217, 234), (203, 216, 234), (202, 213, 232), (211, 223, 238), (196, 208, 222), (195, 208, 223), (204, 220, 233), (205, 223, 233), (203, 222, 229), (207, 227, 233), (207, 226, 233), (211, 226, 238), (212, 225, 239), (215, 226, 239), (217, 225, 237), (219, 224, 235), (220, 224, 234), (221, 223, 234), (221, 224, 234), (220, 226, 234), (219, 226, 234), (219, 226, 234), (220, 227, 234), (220, 227, 233), (221, 227, 233), (221, 227, 232), (223, 228, 232), (222, 227, 231), (221, 227, 231), (221, 228, 232), (220, 228, 232), (220, 228, 233), (220, 228, 233), (219, 228, 233), (220, 228, 233), (221, 227, 232), (221, 227, 232), (222, 228, 234), (221, 229, 235), (220, 229, 235), (221, 229, 235), (222, 228, 233), (223, 228, 231), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (191, 200, 217), (189, 201, 223), (187, 204, 220), (186, 205, 219), (188, 206, 221), (189, 205, 221), (192, 206, 223), (194, 207, 223), (192, 207, 220), (193, 207, 220), (195, 206, 223), (198, 207, 225), (199, 206, 226), (200, 207, 227), (199, 207, 226), (199, 209, 226), (198, 211, 225), (198, 213, 224), (197, 214, 222), (198, 215, 222), (200, 216, 223), (202, 216, 225), (203, 216, 226), (205, 216, 227), (207, 218, 228), (206, 216, 226), (207, 218, 228), (204, 215, 225), (199, 211, 222), (205, 217, 228), (211, 223, 235), (207, 220, 231), (206, 220, 231), (208, 222, 234), (211, 224, 238), (207, 220, 234), (208, 221, 236), (213, 225, 240), (209, 220, 234), (204, 215, 228), (206, 217, 226), (216, 228, 234), (203, 216, 223), (207, 222, 229), (203, 219, 225), (213, 230, 236), (214, 232, 237), (204, 222, 227), (210, 227, 236), (213, 227, 237), (214, 227, 235), (216, 226, 234), (217, 226, 232), (218, 226, 231), (219, 225, 231), (219, 225, 232), (220, 226, 233), (219, 226, 234), (219, 226, 233), (219, 226, 232), (219, 226, 232), (221, 227, 233), (221, 227, 232), (222, 227, 231), (222, 227, 231), (221, 227, 232), (221, 227, 232), (220, 228, 233), (220, 227, 233), (220, 228, 233), (219, 228, 233), (220, 228, 233), (221, 227, 232), (221, 227, 232), (221, 227, 233), (220, 228, 234), (220, 229, 235), (221, 229, 235), (222, 228, 233), (223, 228, 231), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (191, 200, 217), (189, 201, 223), (186, 203, 219), (186, 205, 219), (187, 205, 220), (189, 205, 221), (192, 206, 223), (194, 207, 223), (193, 206, 220), (194, 206, 220), (196, 206, 223), (196, 206, 225), (198, 206, 226), (199, 207, 227), (198, 208, 226), (197, 208, 225), (199, 211, 224), (198, 212, 222), (198, 214, 221), (199, 215, 221), (201, 216, 223), (201, 215, 224), (203, 216, 227), (203, 215, 227), (205, 216, 225), (204, 215, 223), (208, 219, 228), (210, 221, 231), (208, 219, 231), (209, 220, 233), (210, 220, 235), (206, 216, 231), (207, 217, 232), (208, 218, 233), (211, 221, 236), (211, 222, 235), (211, 223, 236), (211, 223, 236), (208, 220, 232), (207, 220, 229), (207, 222, 227), (208, 223, 226), (197, 212, 216), (209, 224, 229), (207, 222, 227), (208, 223, 228), (206, 221, 226), (213, 228, 233), (212, 227, 232), (213, 226, 232), (215, 227, 231), (216, 227, 230), (217, 227, 229), (217, 226, 229), (218, 226, 230), (218, 226, 231), (218, 226, 232), (218, 225, 232), (218, 226, 232), (219, 227, 232), (219, 227, 232), (220, 226, 232), (220, 226, 231), (220, 226, 231), (220, 226, 231), (220, 226, 231), (220, 226, 232), (219, 226, 232), (219, 226, 232), (219, 227, 233), (218, 227, 233), (219, 227, 232), (221, 227, 232), (221, 227, 232), (221, 227, 233), (220, 228, 234), (219, 228, 234), (220, 228, 234), (221, 227, 232), (222, 227, 230), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (191, 200, 217), (188, 200, 222), (186, 203, 219), (185, 204, 218), (186, 204, 219), (188, 204, 220), (191, 205, 222), (193, 206, 223), (194, 206, 221), (194, 206, 221), (195, 206, 224), (195, 206, 225), (196, 207, 226), (197, 208, 226), (197, 209, 226), (197, 209, 224), (199, 211, 223), (199, 212, 222), (199, 212, 221), (199, 213, 222), (200, 214, 224), (201, 215, 226), (201, 214, 228), (202, 216, 228), (205, 219, 228), (203, 217, 225), (203, 217, 227), (205, 217, 229), (206, 217, 231), (208, 217, 233), (210, 217, 234), (211, 217, 234), (212, 218, 234), (212, 218, 234), (210, 216, 231), (210, 218, 231), (207, 218, 230), (205, 219, 229), (207, 223, 232), (208, 225, 233), (206, 226, 232), (203, 224, 229), (201, 220, 226), (203, 219, 226), (207, 220, 228), (208, 219, 228), (203, 213, 220), (215, 224, 228), (216, 226, 227), (217, 226, 226), (216, 226, 225), (216, 226, 226), (216, 226, 227), (217, 227, 229), (216, 227, 230), (217, 226, 231), (217, 226, 232), (217, 226, 232), (217, 226, 232), (218, 226, 231), (218, 226, 231), (218, 225, 231), (219, 225, 231), (219, 225, 231), (220, 226, 232), (220, 226, 232), (219, 226, 232), (219, 226, 232), (219, 226, 233), (219, 226, 233), (218, 227, 233), (219, 227, 233), (221, 227, 232), (221, 227, 232), (221, 227, 233), (220, 228, 234), (219, 228, 234), (220, 228, 234), (221, 227, 232), (222, 227, 230), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (189, 198, 215), (187, 199, 221), (185, 202, 218), (185, 204, 218), (186, 204, 219), (188, 204, 220), (190, 204, 221), (192, 205, 222), (194, 205, 223), (194, 205, 223), (194, 206, 223), (194, 207, 224), (194, 208, 224), (194, 209, 224), (195, 210, 224), (196, 210, 223), (198, 211, 222), (199, 211, 223), (199, 211, 223), (200, 212, 225), (200, 213, 227), (200, 214, 228), (200, 214, 230), (200, 215, 229), (204, 219, 231), (203, 218, 229), (202, 217, 229), (203, 216, 230), (206, 218, 233), (207, 217, 233), (209, 218, 234), (211, 218, 234), (212, 218, 232), (213, 219, 233), (212, 219, 231), (214, 222, 234), (212, 223, 234), (206, 220, 230), (208, 224, 234), (206, 224, 234), (204, 224, 231), (210, 230, 237), (216, 233, 241), (198, 212, 222), (207, 218, 230), (219, 227, 239), (214, 222, 232), (213, 221, 227), (216, 224, 226), (216, 225, 224), (216, 225, 223), (215, 225, 225), (216, 226, 228), (216, 225, 230), (216, 226, 233), (216, 226, 234), (217, 226, 233), (217, 226, 232), (217, 226, 232), (217, 226, 231), (218, 226, 231), (218, 226, 231), (218, 226, 231), (218, 225, 231), (219, 226, 232), (219, 226, 232), (219, 226, 232), (219, 226, 233), (219, 226, 233), (219, 226, 234), (218, 227, 234), (219, 227, 233), (221, 227, 232), (221, 227, 232), (220, 226, 232), (219, 227, 233), (218, 227, 233), (219, 227, 233), (220, 226, 231), (221, 226, 229), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (188, 197, 214), (186, 198, 220), (185, 202, 218), (184, 203, 217), (186, 204, 219), (187, 203, 219), (189, 203, 220), (191, 204, 222), (194, 204, 223), (193, 204, 223), (193, 206, 223), (191, 207, 221), (191, 209, 221), (192, 210, 221), (192, 210, 221), (195, 210, 222), (197, 211, 223), (198, 210, 224), (200, 210, 226), (201, 211, 228), (199, 212, 229), (199, 213, 231), (199, 215, 232), (199, 215, 232), (200, 214, 232), (203, 217, 235), (204, 218, 236), (204, 218, 235), (206, 220, 236), (206, 219, 234), (205, 217, 230), (206, 217, 228), (209, 219, 227), (212, 221, 229), (206, 216, 224), (209, 219, 228), (208, 219, 230), (204, 216, 229), (209, 223, 237), (208, 222, 235), (212, 225, 234), (210, 223, 230), (212, 223, 233), (212, 221, 234), (218, 225, 241), (214, 221, 238), (215, 223, 238), (217, 227, 238), (214, 225, 230), (213, 225, 227), (213, 226, 226), (214, 225, 228), (215, 224, 232), (216, 224, 236), (218, 224, 239), (217, 225, 239), (216, 226, 235), (216, 226, 232), (217, 226, 232), (217, 226, 231), (217, 226, 231), (218, 226, 231), (218, 226, 231), (218, 225, 231), (218, 225, 231), (218, 225, 231), (218, 225, 231), (218, 225, 232), (218, 225, 232), (218, 225, 233), (217, 225, 234), (218, 225, 233), (220, 226, 232), (220, 226, 231), (220, 226, 232), (219, 227, 233), (218, 227, 233), (219, 227, 233), (220, 226, 231), (221, 226, 229), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 1, 0), (0, 0, 0), (1, 0, 1), (2, 0, 2), (2, 0, 2), (1, 0, 0), (0, 1, 0), (0, 2, 4), (188, 197, 214), (186, 198, 220), (184, 201, 217), (184, 203, 217), (186, 204, 219), (187, 203, 219), (189, 203, 220), (190, 202, 221), (194, 204, 224), (194, 204, 223), (191, 205, 222), (191, 208, 221), (190, 210, 220), (190, 210, 219), (192, 211, 220), (193, 210, 221), (197, 211, 223), (199, 210, 225), (200, 210, 228), (200, 210, 229), (199, 211, 231), (199, 213, 232), (199, 215, 233), (199, 215, 234), (198, 212, 233), (202, 215, 237), (202, 216, 236), (199, 214, 232), (201, 217, 233), (202, 217, 230), (201, 216, 227), (203, 217, 225), (205, 217, 222), (210, 221, 226), (207, 218, 223), (211, 222, 230), (212, 223, 234), (207, 219, 233), (209, 222, 238), (206, 218, 233), (210, 220, 230), (215, 224, 232), (211, 219, 230), (216, 224, 237), (218, 224, 242), (213, 219, 238), (215, 223, 241), (211, 222, 235), (213, 225, 232), (212, 226, 229), (212, 226, 228), (213, 225, 230), (214, 224, 234), (216, 223, 239), (218, 224, 242), (218, 224, 241), (216, 226, 236), (216, 226, 232), (217, 226, 232), (217, 226, 231), (217, 226, 231), (217, 226, 231), (218, 226, 231), (218, 225, 231), (218, 225, 231), (218, 225, 231), (218, 225, 231), (218, 225, 232), (218, 225, 232), (218, 225, 233), (217, 225, 234), (218, 225, 233), (220, 226, 232), (220, 226, 231), (220, 226, 232), (219, 227, 233), (218, 227, 233), (219, 227, 233), (219, 225, 230), (220, 225, 228), (0, 1, 3), (0, 0, 1), (1, 0, 0), (1, 0, 0), (1, 0, 0), (1, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0), (0, 0, 0)
);


end package pmod_lcd_pkg;
-------------------------------------------------------------------------------
package body pmod_lcd_pkg is

end package body pmod_lcd_pkg;