library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-------------------------------------------------------------------------------
package pmod_lcd_pkg is

  -- factor for the clock divider , to reduce the SPI clock from the system clock
  constant c_clk_reduce             : integer := 3;
  -- proper reset time
  -- 1 clk = 20 ns ==> 1 us = 50x
  constant c_clk_per_us             : integer :=     50 ; -- clock cycles for 1 us
  constant c_rst_time_act           : integer :=      20 * c_clk_per_us ; -- $9.17   minimum      10 us
  constant c_rst_time_hld           : integer := 125_000 * c_clk_per_us ; -- $9.17   minimum 120_000 us
  constant c_sleep_out              : integer := 125_000 * c_clk_per_us ; -- $9.19.2 minimum 120_000 us

  -- constants found in the LCD controller datasheet
  constant c_bits_565         : integer := 5+6+5;
  constant c_bits_666         : integer := 8+8+8;
  constant c_bits             : integer := c_bits_666;

  -- memory area
  -- the memory is X:132 x Y:162
  constant c_hori             : integer :=  160      ; --! display X
  constant c_vert             : integer :=  132 -26  ; --! display Y
  constant c_ras_xs           : integer :=  1   ;                    --! RAS Xstart
  constant c_ras_xe           : integer :=  c_ras_xs +  c_hori - 1;  --! RAS Xend
  constant c_cas_ys           : integer :=  26  ;                    --! CAS Ystart
  constant c_cas_ye           : integer :=  c_cas_ys +  c_vert - 1;  --! CAS Yend
  constant c_pixl             : integer :=  c_hori * c_vert;         --! total amount of pixels

  -- display area
  constant c_res_x            : integer :=  160      ; --! img X resolution
  constant c_res_y            : integer :=   80      ; --! img Y resolution
  constant c_pixl_img         : integer :=  c_res_x * c_res_y;         --! total amount of pixels

  constant c_SLPOUT           : std_logic_vector(7 downto 0) := x"11";  --! sleep out
  constant c_DISPINV          : std_logic_vector(7 downto 0) := x"21";  --! display inversion
  constant c_DISPOFF          : std_logic_vector(7 downto 0) := x"28";  --! display off
  constant c_DISPON           : std_logic_vector(7 downto 0) := x"29";  --! display on
  constant c_CASET            : std_logic_vector(7 downto 0) := x"2A";  --! column address set
  constant c_RASET            : std_logic_vector(7 downto 0) := x"2B";  --! row address set
  constant c_RAMWR            : std_logic_vector(7 downto 0) := x"2C";  --! RAM write
  constant c_MADCTL           : std_logic_vector(7 downto 0) := x"36";  --! axis control
  constant c_COLMOD           : std_logic_vector(7 downto 0) := x"3A";  --! color mode
  constant c_INVCTR           : std_logic_vector(7 downto 0) := x"B4";  --! display inversion

  -- set display as a landscape mode , and reverse RGB<>BGR
  constant c_MADCTL_P0        : std_logic_vector(7 downto 0) := x"78";  --! parameter 0
  -- set swap dot <> column
  constant c_INVCTR_P0        : std_logic_vector(7 downto 0) := x"03";  --! parameter 0

  -- pre coded RGB values
  constant c_r_color       : std_logic_vector(24-1 downto 0) :=  "11111111" & "00000000" & "00000000" ;
  constant c_g_color       : std_logic_vector(24-1 downto 0) :=  "00000000" & "11111111" & "00000000" ;
  constant c_b_color       : std_logic_vector(24-1 downto 0) :=  "00000000" & "00000000" & "11111111" ;

  -- create arrays for pixel map stores
  type t_raw_arr  is array (integer range <>) of std_logic_vector(24-1 downto 0);     -- raw pixel map
  type t_rgb_arr  is array (integer range <>) of integer range 0 to 255;              -- rgb array
  type t_clr_arr  is array (integer range <>) of t_rgb_arr( 0 to 2);                  -- color array
  type t_cnt_arr  is array (integer range <>) of integer range 0 to c_bits-1;         -- counter array

  constant c_test_map : t_clr_arr( 0 to c_pixl_img-1) :=
  (others => (255, 11, 255));


  constant c_color_map : t_clr_arr( 0 to c_pixl_img-1) :=
((7, 73, 170), (11, 73, 168), (28, 72, 161), (31, 64, 157), (94, 77, 152), (237, 142, 129), (254, 134, 73), (251, 126, 65), (249, 133, 71), (251, 140, 78), (255, 158, 106), (238, 97, 130), (240, 2, 135), (241, 1, 146), (240, 2, 130), (239, 2, 115), (237, 0, 98), (237, 2, 76), (231, 2, 61), (214, 3, 12), (210, 1, 0), (203, 28, 4), (227, 109, 15), (244, 175, 18), (253, 209, 6), (255, 224, 1), (255, 221, 1), (255, 217, 0), (254, 214, 2), (253, 211, 2), (252, 209, 1), (251, 208, 1), (253, 206, 0), (253, 205, 0), (253, 207, 0), (254, 208, 2), (255, 206, 2), (253, 198, 4), (253, 184, 11), (245, 138, 6), (232, 99, 1), (232, 97, 0), (236, 99, 0), (238, 101, 0), (246, 109, 3), (249, 114, 2), (253, 120, 3), (245, 105, 6), (250, 116, 6), (253, 132, 8), (250, 140, 18), (253, 140, 21), (252, 111, 5), (253, 105, 1), (253, 109, 2), (254, 112, 3), (254, 113, 2), (253, 112, 0), (252, 110, 1), (248, 110, 3), (232, 115, 0), (229, 118, 2), (230, 112, 3), (224, 100, 2), (225, 106, 0), (222, 136, 64), (193, 149, 172), (175, 136, 169), (168, 126, 166), (160, 123, 161), (157, 119, 161), (154, 113, 161), (152, 107, 159), (149, 101, 155), (146, 98, 153), (144, 96, 151), (143, 93, 148), (137, 81, 135), (134, 78, 131), (132, 78, 126), (137, 87, 124), (71, 44, 56), (27, 9, 11), (31, 11, 16), (30, 14, 18), (31, 13, 15), (53, 15, 19), (85, 23, 35), (88, 21, 37), (75, 11, 23), (87, 25, 9), (146, 86, 35), (184, 147, 103), (237, 223, 199), (255, 245, 225), (254, 243, 228), (253, 244, 232), (252, 242, 230), (254, 239, 223), (255, 238, 219), (254, 237, 216), (252, 236, 212), (253, 236, 214), (254, 235, 211), (254, 234, 206), (255, 234, 210), (254, 236, 211), (252, 236, 209), (253, 235, 209), (255, 235, 213), (252, 233, 209), (254, 234, 211), (254, 235, 212), (253, 234, 212), (254, 236, 214), (254, 234, 217), (253, 234, 214), (253, 235, 209), (250, 224, 198), (227, 161, 135), (208, 82, 48), (200, 17, 3), (201, 0, 0), (204, 0, 0), (205, 1, 2), (203, 2, 1), (202, 0, 0), (198, 0, 0), (222, 54, 43), (232, 99, 79), (252, 134, 118), (255, 136, 121), (252, 128, 108), (233, 89, 72), (208, 35, 29), (197, 1, 3), (225, 29, 15), (217, 14, 3), (210, 1, 1), (209, 0, 0), (207, 0, 0), (208, 0, 0), (207, 1, 0), (210, 1, 1), (212, 1, 1), (214, 1, 0), (221, 8, 0), (208, 91, 8), (186, 154, 27), (220, 154, 79), (251, 176, 133), (255, 168, 139), (255, 160, 138), (253, 161, 135), (253, 169, 132), (252, 181, 91), (251, 198, 27), (243, 193, 5), (231, 175, 5), (231, 169, 4), (30, 72, 163), (18, 66, 157), (14, 56, 148), (27, 49, 139), (153, 78, 101), (255, 96, 26), (249, 83, 6), (253, 91, 8), (253, 98, 8), (254, 104, 11), (254, 114, 15), (254, 123, 52), (239, 42, 100), (244, 0, 126), (238, 1, 116), (236, 0, 101), (236, 0, 89), (234, 1, 76), (229, 1, 50), (212, 1, 2), (214, 16, 2), (213, 21, 3), (211, 12, 1), (208, 18, 16), (208, 49, 42), (225, 102, 34), (237, 149, 30), (244, 179, 15), (251, 198, 4), (254, 204, 6), (255, 205, 10), (255, 203, 10), (255, 202, 8), (254, 197, 7), (249, 182, 8), (240, 159, 10), (230, 133, 10), (244, 129, 7), (240, 107, 5), (239, 95, 2), (233, 96, 2), (230, 93, 0), (228, 91, 0), (231, 94, 0), (237, 97, 3), (236, 97, 1), (237, 96, 0), (243, 102, 2), (245, 106, 1), (246, 106, 2), (248, 111, 0), (250, 116, 1), (251, 113, 6), (250, 104, 4), (255, 109, 5), (255, 111, 2), (255, 112, 2), (253, 111, 1), (250, 112, 1), (247, 115, 4), (229, 104, 6), (217, 97, 6), (230, 112, 4), (239, 130, 6), (240, 135, 16), (192, 119, 101), (158, 106, 140), (142, 95, 121), (136, 92, 120), (133, 89, 120), (128, 83, 120), (124, 78, 122), (124, 72, 122), (126, 71, 122), (124, 72, 122), (125, 77, 123), (133, 85, 129), (123, 73, 113), (117, 67, 103), (115, 65, 98), (118, 70, 102), (99, 65, 83), (33, 14, 18), (32, 12, 15), (33, 14, 15), (49, 17, 19), (74, 22, 29), (73, 13, 25), (82, 17, 30), (131, 81, 86), (199, 181, 174), (250, 244, 230), (255, 253, 239), (255, 243, 226), (252, 236, 219), (254, 238, 223), (254, 238, 223), (253, 234, 216), (254, 233, 210), (254, 230, 205), (252, 229, 204), (251, 229, 203), (253, 229, 204), (253, 228, 199), (252, 226, 193), (251, 226, 196), (252, 228, 199), (251, 228, 198), (251, 227, 198), (253, 230, 201), (253, 230, 203), (254, 231, 207), (253, 231, 207), (251, 229, 203), (255, 233, 210), (254, 232, 207), (254, 232, 214), (253, 231, 210), (249, 232, 207), (254, 242, 216), (252, 239, 206), (237, 195, 166), (217, 97, 81), (200, 11, 10), (200, 0, 0), (205, 0, 0), (196, 3, 1), (222, 73, 57), (251, 117, 94), (246, 108, 83), (242, 92, 65), (241, 86, 60), (240, 86, 61), (247, 96, 70), (251, 98, 73), (234, 56, 41), (217, 12, 5), (206, 1, 0), (207, 0, 1), (208, 1, 0), (207, 0, 0), (207, 0, 0), (206, 1, 0), (208, 1, 0), (211, 1, 1), (216, 0, 0), (217, 4, 1), (202, 82, 61), (237, 137, 121), (255, 134, 125), (245, 113, 101), (242, 103, 88), (244, 103, 86), (245, 105, 91), (246, 111, 99), (250, 121, 116), (255, 144, 108), (246, 176, 31), (232, 170, 0), (226, 156, 3), (28, 65, 158), (48, 69, 153), (108, 103, 179), (139, 110, 185), (193, 88, 110), (247, 67, 1), (250, 69, 0), (250, 78, 3), (250, 84, 0), (251, 89, 0), (253, 92, 0), (254, 99, 2), (248, 63, 48), (240, 0, 96), (233, 0, 102), (232, 5, 96), (231, 0, 83), (229, 0, 66), (221, 0, 30), (207, 2, 1), (210, 28, 4), (207, 38, 2), (210, 38, 0), (214, 35, 17), (202, 0, 64), (199, 0, 70), (198, 0, 65), (200, 15, 56), (209, 47, 21), (207, 73, 6), (209, 77, 8), (210, 75, 7), (207, 59, 6), (202, 43, 6), (198, 25, 6), (190, 4, 7), (199, 21, 9), (244, 91, 8), (239, 90, 1), (237, 92, 2), (233, 93, 4), (226, 86, 2), (229, 98, 4), (241, 124, 9), (245, 131, 11), (242, 128, 10), (231, 102, 4), (231, 86, 3), (238, 93, 2), (239, 94, 2), (241, 94, 2), (241, 97, 2), (241, 100, 3), (237, 91, 2), (243, 94, 3), (252, 104, 5), (253, 108, 4), (252, 112, 4), (246, 113, 0), (253, 127, 7), (217, 86, 9), (204, 78, 7), (234, 125, 7), (248, 155, 1), (237, 149, 32), (166, 92, 99), (138, 77, 102), (124, 71, 91), (117, 68, 91), (113, 65, 89), (108, 63, 88), (107, 60, 89), (108, 59, 91), (110, 58, 91), (109, 59, 91), (109, 61, 94), (112, 65, 99), (111, 64, 96), (108, 61, 91), (106, 59, 87), (107, 59, 85), (109, 63, 84), (49, 20, 30), (27, 7, 9), (42, 15, 18), (69, 19, 24), (76, 11, 19), (120, 77, 76), (208, 187, 178), (255, 252, 238), (255, 255, 241), (255, 242, 230), (255, 238, 223), (254, 236, 217), (254, 234, 215), (255, 235, 213), (254, 232, 206), (253, 228, 199), (254, 226, 194), (252, 225, 189), (253, 225, 190), (251, 225, 190), (252, 226, 191), (253, 223, 184), (250, 221, 178), (250, 221, 179), (253, 225, 185), (252, 224, 185), (252, 222, 186), (254, 225, 194), (252, 224, 195), (254, 227, 199), (253, 226, 199), (252, 225, 197), (253, 227, 194), (251, 226, 195), (254, 229, 206), (254, 227, 197), (252, 226, 193), (254, 230, 202), (254, 230, 205), (254, 236, 208), (255, 243, 209), (242, 196, 166), (211, 87, 71), (192, 0, 0), (217, 42, 33), (239, 99, 69), (230, 66, 30), (227, 55, 17), (224, 52, 15), (223, 50, 15), (221, 48, 12), (222, 49, 12), (225, 50, 14), (227, 41, 19), (210, 5, 3), (204, 0, 0), (204, 0, 0), (206, 1, 0), (207, 0, 0), (207, 0, 0), (206, 0, 0), (208, 1, 0), (213, 1, 2), (210, 0, 0), (224, 56, 42), (255, 132, 108), (249, 102, 81), (239, 78, 55), (234, 70, 49), (230, 69, 48), (229, 71, 52), (232, 72, 56), (233, 77, 59), (238, 83, 68), (243, 93, 79), (244, 124, 80), (233, 151, 27), (226, 153, 0), (71, 68, 158), (216, 140, 206), (255, 153, 211), (255, 150, 215), (253, 149, 214), (247, 109, 137), (245, 63, 20), (250, 69, 0), (248, 75, 1), (247, 78, 3), (251, 80, 4), (252, 85, 0), (248, 60, 17), (235, 37, 94), (240, 95, 135), (242, 104, 134), (243, 87, 121), (229, 44, 75), (199, 2, 5), (204, 0, 1), (203, 15, 2), (203, 31, 1), (207, 37, 1), (212, 36, 12), (196, 8, 34), (197, 1, 71), (203, 0, 82), (206, 0, 84), (200, 4, 39), (194, 21, 0), (190, 18, 0), (188, 12, 0), (186, 0, 0), (191, 0, 0), (192, 0, 0), (191, 0, 3), (199, 14, 6), (242, 90, 10), (236, 90, 1), (232, 85, 0), (229, 90, 4), (235, 102, 7), (255, 134, 8), (255, 145, 6), (255, 148, 10), (255, 156, 8), (255, 160, 9), (241, 121, 6), (230, 84, 1), (232, 82, 0), (231, 82, 0), (231, 86, 1), (234, 90, 2), (231, 81, 1), (227, 73, 0), (230, 78, 1), (236, 91, 1), (251, 115, 11), (238, 107, 3), (236, 108, 1), (224, 95, 6), (216, 94, 4), (228, 115, 1), (240, 134, 0), (212, 119, 29), (143, 69, 78), (121, 60, 76), (113, 55, 72), (107, 53, 72), (102, 52, 72), (100, 51, 73), (100, 51, 75), (100, 51, 76), (99, 51, 75), (98, 52, 75), (99, 51, 78), (100, 51, 80), (104, 52, 74), (105, 51, 69), (106, 51, 69), (109, 53, 71), (111, 56, 71), (66, 27, 35), (29, 6, 9), (32, 0, 0), (95, 48, 48), (190, 162, 158), (255, 246, 234), (255, 255, 240), (255, 241, 227), (252, 233, 218), (253, 231, 211), (254, 230, 209), (254, 230, 206), (254, 228, 203), (254, 227, 199), (252, 224, 189), (252, 221, 183), (254, 219, 179), (253, 216, 176), (254, 216, 175), (253, 217, 175), (254, 218, 176), (253, 214, 170), (252, 210, 163), (255, 213, 170), (255, 216, 180), (254, 217, 184), (253, 217, 182), (255, 220, 184), (252, 218, 179), (253, 221, 182), (252, 221, 184), (252, 221, 187), (254, 223, 192), (252, 221, 194), (252, 223, 194), (250, 220, 186), (255, 226, 195), (253, 227, 199), (254, 229, 199), (251, 222, 192), (254, 227, 196), (253, 236, 202), (255, 237, 201), (230, 175, 151), (220, 100, 73), (217, 39, 0), (210, 37, 0), (208, 30, 0), (207, 24, 2), (209, 21, 3), (210, 18, 0), (209, 14, 0), (208, 8, 0), (201, 0, 0), (199, 0, 0), (203, 2, 2), (204, 1, 1), (206, 0, 0), (207, 0, 0), (207, 0, 0), (207, 0, 0), (209, 1, 0), (205, 0, 0), (208, 18, 13), (245, 102, 82), (239, 86, 61), (230, 61, 28), (226, 54, 15), (219, 50, 12), (215, 49, 13), (214, 51, 17), (217, 52, 22), (222, 59, 28), (225, 65, 35), (230, 72, 44), (237, 88, 65), (239, 128, 52), (227, 146, 2), (175, 74, 172), (255, 63, 180), (248, 30, 162), (250, 35, 176), (252, 57, 189), (253, 77, 207), (248, 62, 120), (249, 58, 3), (251, 69, 0), (246, 69, 0), (247, 69, 0), (252, 69, 0), (248, 63, 23), (237, 94, 101), (233, 109, 111), (233, 104, 107), (236, 105, 107), (242, 106, 105), (219, 53, 52), (195, 0, 1), (195, 0, 0), (194, 9, 0), (201, 16, 6), (193, 13, 7), (168, 1, 0), (172, 2, 14), (182, 4, 32), (185, 3, 36), (184, 5, 17), (192, 18, 3), (193, 19, 1), (191, 13, 1), (190, 2, 1), (191, 1, 1), (190, 1, 1), (188, 1, 3), (183, 0, 1), (216, 51, 5), (236, 94, 3), (228, 89, 2), (226, 95, 3), (243, 121, 6), (246, 125, 1), (244, 122, 0), (247, 125, 0), (252, 133, 0), (253, 144, 2), (255, 150, 11), (238, 102, 6), (230, 77, 0), (231, 80, 0), (230, 83, 0), (231, 84, 0), (228, 79, 0), (229, 78, 1), (228, 81, 0), (229, 88, 0), (235, 100, 4), (228, 97, 1), (226, 93, 2), (218, 87, 3), (218, 93, 3), (224, 102, 0), (222, 111, 0), (191, 94, 20), (127, 58, 57), (113, 53, 52), (105, 44, 57), (100, 43, 56), (96, 44, 56), (96, 42, 58), (97, 42, 60), (96, 42, 60), (96, 41, 60), (99, 45, 63), (98, 43, 61), (97, 42, 59), (100, 43, 57), (100, 42, 54), (102, 46, 53), (107, 51, 55), (113, 55, 61), (65, 23, 26), (23, 1, 1), (124, 99, 91), (239, 226, 212), (255, 255, 244), (255, 241, 225), (252, 237, 217), (251, 235, 212), (253, 228, 202), (251, 223, 187), (252, 222, 193), (251, 220, 187), (252, 219, 185), (254, 218, 184), (252, 213, 169), (252, 212, 166), (253, 209, 160), (253, 207, 158), (251, 208, 153), (252, 208, 153), (254, 207, 155), (253, 204, 152), (251, 203, 152), (251, 204, 153), (254, 207, 162), (252, 207, 166), (252, 209, 167), (255, 214, 171), (251, 210, 167), (253, 214, 174), (254, 216, 178), (253, 214, 176), (255, 218, 180), (255, 218, 183), (254, 220, 186), (252, 217, 182), (254, 220, 188), (254, 223, 191), (254, 223, 186), (251, 220, 183), (251, 225, 193), (250, 224, 196), (253, 224, 196), (255, 239, 209), (247, 228, 189), (217, 126, 88), (191, 15, 0), (199, 3, 0), (198, 3, 1), (198, 2, 1), (196, 2, 0), (198, 1, 0), (197, 0, 1), (193, 1, 2), (189, 3, 2), (193, 3, 3), (203, 1, 4), (209, 0, 1), (209, 0, 0), (208, 0, 0), (208, 0, 0), (208, 0, 0), (207, 12, 8), (224, 64, 48), (239, 82, 55), (225, 52, 14), (216, 41, 5), (211, 33, 2), (205, 28, 0), (202, 28, 0), (204, 30, 0), (205, 34, 2), (207, 41, 5), (213, 47, 10), (217, 52, 15), (225, 61, 26), (237, 99, 39), (231, 141, 7), (228, 100, 168), (245, 0, 158), (250, 0, 170), (251, 0, 170), (252, 0, 170), (249, 0, 165), (249, 13, 156), (251, 38, 33), (246, 62, 3), (245, 94, 49), (245, 113, 59), (241, 82, 34), (220, 36, 21), (221, 61, 63), (223, 66, 65), (222, 68, 63), (222, 70, 62), (224, 76, 64), (232, 75, 63), (199, 20, 17), (180, 0, 0), (181, 1, 1), (179, 1, 2), (172, 0, 1), (166, 2, 0), (166, 1, 0), (168, 2, 0), (170, 1, 0), (172, 1, 0), (184, 11, 3), (190, 12, 3), (188, 4, 0), (190, 1, 2), (188, 0, 3), (187, 0, 0), (186, 1, 1), (181, 0, 4), (203, 47, 14), (228, 104, 6), (217, 91, 1), (222, 96, 3), (236, 115, 4), (232, 109, 1), (230, 105, 0), (234, 107, 1), (243, 112, 1), (249, 120, 1), (254, 134, 6), (248, 116, 8), (225, 73, 2), (229, 76, 5), (228, 77, 3), (226, 75, 0), (227, 77, 0), (228, 80, 0), (228, 83, 1), (226, 86, 1), (224, 87, 0), (221, 85, 3), (221, 83, 6), (204, 64, 4), (213, 88, 1), (209, 104, 30), (209, 119, 108), (172, 95, 90), (116, 44, 39), (111, 46, 44), (104, 43, 49), (99, 41, 50), (96, 40, 50), (96, 39, 51), (97, 38, 51), (97, 37, 51), (100, 38, 52), (103, 41, 55), (98, 37, 48), (100, 41, 48), (101, 44, 49), (100, 44, 47), (101, 46, 44), (106, 50, 45), (99, 40, 37), (79, 38, 31), (173, 156, 143), (255, 249, 235), (255, 244, 227), (253, 233, 215), (253, 232, 213), (254, 229, 212), (253, 224, 201), (251, 214, 177), (249, 209, 160), (254, 213, 175), (252, 210, 170), (254, 209, 165), (255, 207, 165), (252, 203, 151), (251, 201, 147), (253, 199, 140), (253, 198, 139), (251, 198, 134), (254, 198, 140), (254, 198, 135), (253, 196, 131), (252, 196, 135), (252, 197, 133), (253, 202, 144), (252, 203, 149), (251, 205, 152), (254, 206, 157), (250, 203, 149), (254, 207, 164), (253, 208, 163), (251, 208, 161), (254, 210, 163), (253, 212, 169), (253, 214, 176), (252, 213, 176), (254, 217, 181), (254, 217, 182), (254, 217, 179), (253, 215, 177), (251, 219, 187), (250, 219, 190), (252, 221, 190), (252, 226, 197), (253, 233, 208), (255, 243, 216), (226, 164, 131), (194, 16, 15), (198, 0, 0), (200, 0, 0), (196, 0, 0), (195, 1, 0), (192, 1, 2), (190, 1, 2), (187, 2, 3), (175, 2, 1), (179, 1, 1), (196, 1, 2), (197, 1, 1), (198, 1, 1), (199, 1, 1), (202, 2, 2), (231, 40, 26), (237, 78, 47), (221, 52, 14), (212, 32, 0), (207, 22, 3), (201, 15, 4), (195, 9, 1), (194, 9, 1), (198, 13, 1), (197, 20, 2), (193, 22, 1), (201, 28, 0), (208, 35, 2), (215, 41, 5), (227, 72, 14), (231, 137, 6), (255, 173, 128), (245, 107, 144), (247, 6, 159), (251, 0, 162), (249, 0, 155), (250, 0, 145), (252, 0, 145), (245, 21, 81), (245, 117, 109), (246, 180, 181), (246, 199, 198), (247, 194, 194), (235, 127, 119), (213, 45, 42), (213, 45, 34), (213, 48, 21), (214, 49, 19), (218, 53, 18), (220, 58, 24), (206, 37, 32), (167, 5, 7), (160, 1, 0), (163, 2, 0), (163, 1, 0), (165, 2, 1), (167, 1, 0), (167, 2, 0), (170, 1, 2), (169, 0, 2), (209, 45, 13), (210, 46, 9), (181, 0, 0), (186, 1, 1), (187, 0, 1), (186, 0, 1), (180, 0, 2), (192, 26, 10), (226, 102, 13), (216, 99, 1), (215, 89, 1), (223, 97, 7), (232, 107, 5), (226, 99, 0), (225, 96, 0), (227, 95, 2), (233, 100, 3), (239, 105, 3), (247, 115, 4), (243, 108, 6), (213, 68, 1), (215, 69, 2), (215, 66, 1), (217, 65, 0), (225, 75, 1), (227, 80, 1), (224, 82, 2), (219, 82, 1), (219, 80, 3), (219, 81, 4), (205, 71, 5), (197, 60, 2), (196, 84, 36), (170, 93, 130), (171, 104, 180), (154, 86, 131), (110, 40, 34), (110, 43, 30), (105, 43, 41), (101, 42, 45), (99, 41, 45), (100, 41, 45), (101, 41, 45), (100, 41, 45), (102, 43, 45), (103, 45, 46), (102, 43, 42), (103, 44, 42), (103, 47, 38), (102, 46, 36), (103, 47, 35), (92, 33, 20), (117, 67, 54), (225, 202, 185), (255, 253, 234), (254, 235, 215), (253, 231, 209), (252, 227, 204), (255, 220, 200), (254, 215, 189), (255, 214, 178), (255, 206, 164), (254, 201, 155), (253, 202, 150), (255, 201, 148), (254, 200, 147), (254, 199, 144), (251, 194, 131), (253, 192, 127), (253, 189, 120), (253, 188, 116), (253, 188, 115), (255, 190, 121), (254, 191, 119), (252, 188, 109), (251, 185, 104), (254, 187, 120), (254, 194, 128), (251, 195, 130), (251, 197, 133), (253, 199, 138), (249, 194, 122), (253, 199, 138), (248, 198, 139), (249, 200, 143), (252, 204, 152), (254, 205, 156), (254, 205, 159), (250, 204, 159), (255, 210, 166), (253, 209, 170), (253, 211, 172), (254, 212, 172), (253, 212, 171), (253, 215, 172), (250, 217, 173), (252, 221, 188), (253, 222, 195), (252, 224, 198), (255, 244, 215), (239, 190, 169), (199, 37, 31), (191, 0, 0), (196, 0, 0), (195, 1, 0), (192, 1, 2), (191, 1, 3), (185, 1, 2), (171, 1, 0), (165, 2, 0), (168, 1, 1), (169, 1, 1), (174, 0, 1), (179, 1, 1), (190, 5, 4), (205, 19, 7), (225, 48, 14), (213, 35, 0), (207, 18, 3), (199, 4, 3), (197, 1, 3), (194, 0, 1), (191, 0, 1), (192, 2, 1), (190, 4, 2), (186, 3, 1), (193, 7, 2), (200, 15, 4), (209, 25, 1), (217, 64, 3), (221, 139, 5), (251, 105, 26), (252, 131, 67), (246, 52, 127), (249, 0, 153), (251, 0, 152), (248, 0, 147), (250, 0, 142), (243, 29, 113), (243, 130, 139), (239, 146, 137), (241, 153, 141), (243, 165, 151), (251, 183, 163), (225, 89, 73), (204, 20, 6), (208, 31, 3), (205, 33, 2), (208, 35, 0), (207, 31, 4), (207, 31, 36), (175, 12, 20), (157, 0, 0), (162, 1, 0), (161, 1, 0), (162, 1, 0), (162, 2, 1), (161, 3, 1), (166, 1, 3), (168, 1, 2), (216, 58, 11), (231, 75, 6), (202, 27, 6), (185, 2, 1), (186, 0, 2), (186, 0, 3), (177, 0, 2), (204, 62, 13), (219, 103, 2), (211, 89, 1), (212, 85, 1), (218, 90, 4), (230, 101, 5), (227, 95, 0), (227, 94, 1), (227, 93, 1), (231, 95, 1), (233, 99, 0), (239, 104, 2), (232, 93, 9), (211, 70, 1), (214, 75, 1), (216, 76, 1), (211, 68, 2), (208, 64, 2), (217, 74, 3), (218, 78, 2), (219, 81, 2), (222, 81, 2), (222, 88, 1), (229, 113, 3), (225, 124, 9), (155, 62, 55), (120, 43, 99), (120, 52, 97), (116, 48, 87), (110, 40, 39), (110, 44, 22), (107, 44, 36), (107, 44, 43), (105, 43, 44), (104, 43, 45), (105, 45, 45), (106, 47, 44), (108, 50, 44), (108, 50, 39), (107, 49, 34), (108, 50, 36), (107, 50, 35), (106, 48, 33), (96, 31, 17), (135, 85, 68), (242, 220, 198), (255, 246, 225), (252, 230, 211), (253, 228, 208), (251, 223, 199), (251, 218, 188), (254, 210, 176), (254, 204, 166), (253, 202, 151), (252, 199, 138), (252, 195, 136), (253, 194, 131), (254, 190, 123), (253, 190, 124), (253, 187, 119), (252, 182, 107), (255, 183, 107), (253, 180, 103), (253, 179, 99), (253, 180, 102), (255, 182, 106), (255, 180, 103), (251, 176, 87), (251, 178, 81), (255, 181, 103), (255, 185, 108), (253, 183, 106), (254, 184, 108), (255, 186, 112), (253, 184, 109), (254, 191, 129), (252, 189, 124), (253, 191, 126), (254, 197, 139), (254, 198, 142), (253, 199, 140), (249, 198, 135), (253, 203, 149), (252, 204, 155), (251, 205, 157), (252, 207, 161), (254, 210, 164), (255, 213, 171), (251, 211, 173), (250, 213, 169), (254, 217, 184), (254, 220, 189), (250, 220, 187), (255, 239, 206), (243, 205, 171), (195, 46, 39), (188, 0, 0), (196, 1, 0), (192, 1, 1), (188, 1, 3), (180, 1, 2), (171, 1, 1), (168, 2, 1), (167, 2, 2), (167, 2, 1), (170, 0, 0), (175, 0, 0), (188, 7, 3), (202, 21, 7), (212, 36, 5), (208, 24, 0), (203, 6, 3), (197, 0, 1), (195, 0, 0), (193, 0, 0), (192, 1, 1), (191, 1, 1), (190, 0, 2), (193, 0, 3), (196, 0, 1), (197, 0, 1), (202, 4, 2), (217, 58, 15), (223, 134, 17), (244, 74, 0), (251, 90, 1), (250, 69, 65), (245, 0, 142), (247, 1, 149), (242, 5, 140), (237, 0, 111), (235, 33, 82), (239, 99, 93), (236, 102, 84), (235, 106, 75), (234, 112, 77), (242, 126, 93), (233, 93, 66), (197, 4, 0), (203, 6, 1), (199, 10, 2), (199, 9, 2), (196, 5, 16), (193, 13, 43), (167, 6, 14), (154, 0, 0), (158, 1, 0), (160, 1, 0), (160, 1, 2), (154, 0, 0), (150, 0, 0), (159, 0, 1), (161, 0, 0), (202, 44, 10), (227, 68, 7), (211, 46, 11), (180, 10, 5), (173, 1, 3), (180, 1, 5), (175, 0, 3), (206, 63, 13), (215, 96, 2), (208, 83, 2), (209, 82, 2), (214, 82, 2), (220, 85, 6), (232, 95, 8), (231, 96, 0), (231, 96, 0), (230, 95, 0), (232, 99, 0), (230, 95, 2), (215, 75, 1), (214, 73, 2), (217, 80, 3), (217, 83, 2), (209, 76, 4), (192, 57, 0), (199, 63, 2), (204, 66, 3), (204, 67, 3), (217, 88, 5), (237, 127, 5), (244, 144, 3), (229, 140, 7), (113, 24, 20), (84, 3, 48), (88, 19, 63), (81, 13, 52), (92, 25, 31), (113, 46, 26), (113, 46, 35), (114, 47, 40), (113, 47, 41), (112, 48, 42), (113, 50, 41), (115, 53, 38), (116, 55, 39), (115, 55, 37), (113, 52, 34), (113, 53, 32), (113, 52, 29), (101, 35, 11), (149, 96, 74), (248, 227, 204), (255, 241, 217), (250, 228, 206), (250, 222, 200), (252, 219, 194), (254, 211, 178), (251, 203, 161), (253, 201, 149), (253, 197, 147), (252, 194, 135), (252, 190, 121), (253, 186, 119), (254, 184, 116), (252, 181, 108), (254, 182, 110), (254, 179, 102), (253, 175, 84), (255, 176, 89), (252, 174, 84), (251, 173, 81), (252, 174, 82), (255, 177, 87), (254, 172, 82), (250, 169, 69), (252, 174, 74), (254, 175, 88), (254, 176, 91), (254, 176, 92), (255, 177, 96), (253, 176, 85), (252, 177, 91), (253, 183, 108), (252, 182, 101), (253, 182, 111), (255, 188, 127), (255, 190, 128), (254, 191, 128), (250, 191, 119), (253, 193, 134), (254, 196, 143), (254, 198, 146), (253, 200, 150), (254, 204, 153), (252, 205, 160), (252, 207, 167), (251, 210, 164), (252, 212, 166), (252, 214, 177), (249, 213, 177), (248, 212, 177), (255, 234, 200), (246, 210, 184), (200, 46, 37), (191, 0, 0), (188, 4, 2), (182, 0, 0), (175, 0, 1), (173, 1, 2), (169, 1, 1), (167, 0, 1), (167, 0, 0), (182, 10, 4), (199, 27, 11), (211, 36, 9), (217, 40, 6), (210, 34, 2), (202, 17, 0), (199, 1, 1), (196, 0, 1), (194, 0, 1), (194, 0, 2), (193, 1, 2), (192, 1, 3), (192, 0, 3), (194, 0, 3), (197, 0, 1), (199, 0, 1), (199, 3, 0), (234, 58, 33), (245, 93, 48), (238, 64, 0), (243, 70, 1), (241, 64, 22), (238, 59, 110), (245, 124, 155), (243, 147, 177), (234, 99, 123), (224, 46, 57), (236, 81, 71), (229, 89, 63), (230, 90, 48), (231, 92, 40), (234, 98, 35), (214, 60, 27), (183, 2, 1), (193, 16, 11), (181, 2, 17), (181, 0, 25), (178, 4, 20), (162, 8, 15), (149, 0, 1), (153, 2, 1), (156, 4, 2), (155, 0, 0), (159, 0, 1), (169, 13, 7), (177, 19, 11), (169, 9, 5), (154, 0, 0), (176, 16, 7), (199, 36, 9), (162, 5, 1), (145, 0, 2), (142, 0, 0), (155, 3, 2), (180, 2, 7), (201, 45, 6), (220, 92, 3), (209, 81, 1), (211, 82, 5), (204, 69, 3), (194, 55, 1), (209, 69, 8), (223, 85, 6), (226, 87, 6), (225, 85, 6), (222, 81, 3), (208, 66, 2), (206, 62, 3), (214, 72, 4), (216, 79, 3), (216, 85, 3), (210, 80, 3), (195, 63, 1), (200, 64, 6), (197, 59, 1), (188, 55, 0), (197, 72, 0), (229, 119, 2), (231, 128, 0), (227, 132, 6), (118, 41, 46), (98, 36, 117), (106, 46, 140), (83, 29, 96), (58, 11, 36), (99, 37, 30), (119, 48, 35), (117, 49, 35), (119, 52, 36), (120, 55, 36), (122, 58, 34), (124, 61, 35), (124, 60, 36), (121, 57, 35), (119, 55, 31), (119, 56, 27), (105, 39, 11), (146, 98, 72), (251, 230, 209), (255, 234, 211), (254, 223, 197), (254, 217, 183), (253, 209, 175), (254, 208, 171), (255, 200, 151), (254, 193, 141), (254, 190, 134), (254, 189, 132), (255, 187, 124), (254, 181, 112), (254, 178, 106), (254, 177, 102), (253, 175, 96), (255, 176, 98), (254, 172, 86), (252, 168, 71), (255, 171, 80), (252, 167, 71), (252, 167, 65), (253, 168, 67), (254, 169, 69), (251, 166, 59), (252, 167, 59), (255, 170, 72), (255, 170, 77), (254, 171, 75), (252, 171, 74), (255, 173, 88), (253, 172, 80), (253, 174, 85), (255, 176, 87), (251, 173, 78), (252, 173, 87), (253, 178, 101), (254, 181, 105), (254, 182, 111), (252, 182, 108), (255, 186, 123), (255, 189, 129), (255, 192, 134), (254, 195, 138), (254, 197, 141), (254, 199, 147), (251, 201, 148), (251, 206, 158), (254, 208, 167), (251, 205, 162), (254, 207, 165), (250, 203, 159), (248, 206, 167), (255, 231, 204), (245, 201, 167), (182, 36, 27), (169, 0, 0), (175, 1, 0), (175, 1, 0), (173, 1, 1), (169, 0, 2), (171, 3, 1), (196, 29, 8), (212, 44, 11), (214, 46, 12), (215, 41, 10), (209, 28, 6), (195, 12, 1), (199, 9, 4), (197, 2, 2), (194, 1, 2), (194, 1, 3), (193, 1, 2), (194, 0, 2), (193, 0, 2), (194, 0, 2), (196, 1, 3), (197, 0, 2), (197, 0, 0), (207, 11, 5), (232, 46, 14), (234, 54, 19), (240, 58, 3), (241, 57, 0), (238, 61, 5), (246, 109, 81), (245, 152, 132), (240, 165, 151), (249, 185, 166), (236, 118, 96), (221, 54, 23), (233, 76, 38), (231, 80, 34), (229, 81, 18), (219, 67, 9), (182, 12, 11), (180, 18, 13), (229, 145, 21), (213, 122, 18), (197, 98, 18), (218, 135, 15), (209, 135, 14), (152, 37, 6), (142, 4, 2), (146, 3, 1), (154, 3, 2), (198, 37, 17), (219, 55, 21), (219, 53, 18), (215, 49, 16), (186, 29, 11), (161, 1, 2), (163, 0, 1), (152, 0, 1), (152, 10, 9), (149, 9, 5), (142, 3, 0), (174, 0, 6), (187, 14, 6), (210, 68, 8), (209, 76, 0), (208, 77, 7), (205, 75, 5), (208, 78, 5), (206, 75, 1), (207, 74, 1), (208, 75, 2), (213, 77, 4), (214, 75, 3), (211, 73, 2), (206, 67, 3), (206, 62, 3), (211, 72, 3), (213, 81, 5), (203, 71, 1), (198, 66, 0), (198, 70, 5), (173, 52, 5), (160, 47, 15), (164, 55, 17), (197, 91, 9), (217, 108, 0), (162, 83, 27), (92, 37, 99), (91, 37, 136), (84, 31, 144), (67, 25, 101), (44, 10, 46), (51, 11, 21), (101, 44, 32), (117, 53, 31), (122, 56, 34), (125, 57, 33), (129, 64, 30), (131, 66, 34), (127, 61, 31), (124, 58, 30), (122, 58, 27), (110, 45, 9), (142, 91, 59), (248, 227, 206), (254, 235, 213), (251, 221, 194), (252, 215, 178), (251, 205, 160), (255, 201, 165), (255, 197, 154), (253, 187, 129), (254, 183, 125), (253, 183, 120), (252, 182, 122), (253, 178, 112), (255, 173, 98), (255, 172, 98), (252, 170, 90), (252, 168, 81), (254, 167, 81), (253, 164, 71), (252, 163, 61), (255, 165, 68), (253, 162, 64), (251, 160, 52), (253, 160, 57), (254, 160, 64), (251, 161, 47), (252, 163, 49), (253, 163, 63), (253, 162, 63), (254, 166, 62), (249, 164, 54), (254, 167, 73), (254, 168, 77), (254, 169, 84), (254, 169, 78), (251, 168, 68), (252, 169, 79), (251, 169, 83), (252, 172, 87), (253, 175, 90), (253, 176, 92), (254, 180, 107), (253, 182, 113), (253, 185, 122), (254, 190, 129), (254, 194, 133), (255, 196, 140), (251, 196, 139), (249, 200, 147), (254, 204, 161), (254, 201, 158), (254, 202, 157), (251, 200, 149), (249, 198, 144), (254, 208, 172), (255, 228, 193), (237, 184, 149), (167, 20, 14), (176, 0, 0), (177, 2, 1), (172, 0, 0), (170, 1, 2), (201, 35, 13), (217, 50, 12), (210, 40, 6), (202, 32, 4), (199, 20, 4), (189, 3, 1), (172, 0, 0), (181, 2, 2), (197, 3, 4), (195, 1, 1), (192, 2, 2), (192, 2, 2), (193, 0, 0), (194, 0, 0), (195, 1, 1), (196, 1, 1), (196, 1, 1), (197, 0, 1), (203, 2, 3), (206, 8, 0), (213, 22, 0), (237, 43, 0), (238, 58, 8), (235, 69, 18), (234, 82, 45), (237, 91, 63), (237, 100, 69), (237, 114, 77), (238, 116, 73), (207, 37, 4), (210, 29, 4), (208, 34, 12), (201, 33, 7), (185, 8, 15), (171, 0, 12), (189, 49, 15), (238, 199, 12), (234, 208, 4), (230, 203, 2), (223, 195, 2), (224, 194, 4), (189, 122, 30), (146, 26, 31), (143, 11, 8), (175, 22, 8), (207, 42, 7), (197, 30, 0), (194, 21, 1), (186, 8, 0), (188, 16, 6), (174, 13, 9), (175, 26, 8), (204, 67, 13), (209, 72, 11), (196, 53, 11), (180, 34, 6), (168, 12, 3), (164, 0, 4), (173, 22, 7), (212, 86, 12), (232, 113, 5), (235, 120, 1), (238, 123, 1), (239, 121, 1), (239, 118, 2), (243, 120, 4), (246, 123, 3), (247, 128, 3), (248, 131, 6), (248, 126, 5), (234, 103, 6), (205, 73, 5), (191, 61, 3), (193, 63, 0), (202, 69, 4), (162, 55, 5), (114, 26, 27), (110, 33, 56), (125, 50, 87), (154, 71, 87), (162, 76, 42), (78, 17, 52), (61, 5, 82), (67, 3, 89), (65, 7, 96), (61, 14, 78), (49, 13, 48), (29, 3, 26), (71, 31, 36), (112, 49, 34), (119, 55, 27), (128, 60, 30), (129, 61, 27), (123, 58, 24), (121, 55, 23), (120, 56, 25), (106, 43, 13), (127, 72, 38), (241, 215, 192), (255, 236, 213), (247, 217, 187), (252, 213, 181), (251, 205, 165), (249, 198, 148), (251, 196, 150), (254, 189, 131), (251, 178, 107), (254, 178, 110), (254, 174, 106), (253, 174, 104), (254, 169, 94), (254, 164, 80), (254, 165, 77), (253, 164, 76), (253, 162, 71), (254, 160, 66), (254, 158, 61), (253, 159, 50), (255, 159, 56), (252, 155, 46), (251, 155, 39), (253, 158, 51), (255, 158, 58), (252, 158, 42), (250, 158, 43), (252, 160, 57), (254, 160, 59), (253, 161, 49), (249, 159, 36), (254, 163, 61), (254, 164, 72), (253, 163, 70), (253, 163, 64), (252, 163, 59), (254, 165, 80), (253, 167, 74), (255, 169, 78), (253, 169, 73), (252, 170, 67), (253, 171, 82), (253, 175, 94), (254, 179, 110), (254, 181, 113), (254, 185, 120), (255, 188, 125), (251, 186, 121), (253, 192, 139), (253, 195, 143), (252, 195, 144), (251, 195, 147), (254, 201, 151), (250, 197, 142), (252, 201, 155), (253, 208, 168), (255, 228, 180), (222, 151, 115), (172, 3, 0), (177, 1, 1), (171, 0, 0), (187, 20, 9), (213, 49, 16), (202, 36, 1), (193, 23, 2), (182, 9, 2), (180, 1, 1), (175, 0, 0), (165, 3, 0), (157, 3, 0), (170, 2, 1), (186, 0, 3), (191, 1, 1), (189, 2, 2), (189, 0, 1), (190, 0, 1), (190, 0, 1), (189, 0, 1), (187, 0, 0), (192, 2, 0), (201, 13, 8), (207, 21, 16), (211, 24, 17), (238, 73, 45), (251, 111, 58), (254, 134, 92), (251, 133, 97), (240, 110, 66), (229, 78, 19), (236, 82, 17), (228, 75, 23), (199, 37, 4), (191, 23, 0), (170, 0, 2), (172, 0, 11), (172, 0, 12), (174, 22, 2), (210, 131, 14), (225, 192, 7), (227, 194, 7), (226, 193, 2), (223, 194, 0), (221, 183, 8), (213, 145, 37), (169, 53, 43), (165, 39, 31), (181, 25, 13), (185, 10, 1), (180, 2, 1), (174, 2, 5), (193, 37, 19), (223, 84, 35), (236, 107, 32), (238, 116, 20), (241, 117, 5), (232, 103, 1), (220, 86, 4), (204, 62, 5), (189, 35, 5), (181, 29, 3), (213, 80, 10), (245, 128, 11), (243, 130, 2), (242, 127, 1), (245, 127, 1), (248, 129, 1), (251, 131, 0), (254, 133, 1), (255, 136, 0), (255, 139, 1), (255, 141, 2), (255, 144, 1), (255, 147, 2), (245, 129, 11), (201, 75, 8), (181, 54, 2), (173, 53, 6), (102, 22, 9), (94, 20, 39), (107, 27, 54), (117, 48, 84), (128, 70, 122), (105, 48, 98), (41, 0, 33), (57, 5, 42), (65, 12, 57), (57, 7, 54), (43, 0, 51), (46, 7, 48), (39, 10, 36), (60, 17, 32), (99, 33, 38), (91, 29, 12), (91, 39, 6), (117, 65, 23), (129, 74, 36), (109, 56, 18), (97, 31, 0), (117, 51, 9), (219, 192, 163), (255, 237, 215), (254, 215, 189), (255, 207, 178), (255, 202, 164), (252, 194, 145), (255, 189, 139), (251, 184, 130), (251, 178, 108), (251, 169, 89), (253, 170, 95), (253, 168, 92), (253, 167, 89), (253, 163, 76), (254, 157, 63), (254, 158, 59), (254, 158, 61), (254, 158, 60), (255, 155, 60), (253, 152, 47), (250, 151, 27), (254, 154, 32), (251, 149, 26), (252, 151, 25), (254, 153, 34), (254, 154, 45), (253, 151, 30), (254, 151, 28), (254, 154, 53), (253, 156, 56), (252, 156, 42), (251, 155, 36), (255, 157, 53), (253, 158, 59), (253, 159, 55), (253, 158, 49), (252, 158, 45), (254, 162, 63), (253, 163, 62), (254, 164, 73), (252, 164, 63), (252, 164, 60), (255, 166, 76), (254, 168, 81), (254, 171, 89), (254, 175, 95), (254, 178, 101), (255, 182, 106), (250, 181, 103), (253, 186, 125), (254, 189, 133), (253, 190, 130), (254, 193, 139), (255, 196, 145), (251, 194, 140), (251, 196, 145), (253, 200, 154), (255, 202, 158), (255, 220, 173), (207, 102, 78), (171, 0, 0), (173, 1, 1), (197, 31, 10), (197, 35, 2), (185, 19, 0), (175, 5, 2), (171, 0, 1), (168, 1, 0), (164, 1, 0), (162, 2, 0), (157, 2, 0), (153, 2, 1), (158, 1, 2), (166, 0, 6), (182, 3, 3), (181, 3, 1), (179, 3, 0), (176, 2, 0), (176, 3, 1), (196, 25, 13), (218, 51, 34), (231, 72, 52), (238, 82, 63), (241, 84, 69), (251, 114, 192), (243, 101, 87), (247, 110, 55), (253, 122, 73), (254, 128, 76), (241, 90, 37), (222, 56, 9), (204, 38, 1), (199, 34, 2), (192, 33, 5), (215, 113, 16), (208, 106, 13), (201, 100, 14), (210, 149, 13), (211, 167, 3), (210, 168, 0), (216, 181, 3), (217, 183, 3), (209, 154, 46), (186, 90, 80), (162, 48, 53), (135, 16, 9), (140, 29, 17), (158, 15, 15), (174, 0, 2), (178, 10, 6), (227, 91, 39), (247, 133, 43), (237, 121, 16), (228, 108, 7), (222, 100, 2), (221, 93, 1), (222, 91, 0), (223, 92, 2), (220, 84, 8), (206, 65, 5), (221, 99, 7), (245, 134, 9), (241, 127, 2), (239, 124, 2), (244, 124, 2), (247, 125, 2), (249, 126, 2), (250, 129, 1), (252, 130, 0), (253, 134, 1), (255, 136, 1), (255, 137, 2), (253, 140, 2), (254, 141, 0), (255, 145, 2), (252, 137, 9), (197, 71, 9), (127, 21, 3), (84, 20, 6), (99, 27, 28), (107, 27, 41), (108, 32, 57), (95, 34, 73), (94, 48, 66), (158, 128, 95), (210, 200, 127), (224, 216, 139), (208, 195, 128), (151, 129, 98), (64, 27, 45), (35, 0, 37), (54, 3, 28), (89, 15, 20), (112, 63, 32), (185, 167, 106), (232, 222, 135), (243, 237, 149), (227, 219, 148), (195, 163, 87), (222, 181, 121), (255, 236, 217), (253, 215, 176), (252, 207, 166), (253, 200, 157), (252, 195, 137), (250, 183, 121), (255, 178, 122), (252, 174, 109), (252, 166, 87), (251, 162, 71), (253, 162, 82), (253, 161, 81), (253, 159, 77), (251, 156, 62), (254, 151, 47), (254, 151, 40), (253, 151, 46), (253, 152, 52), (254, 151, 49), (252, 148, 25), (250, 145, 3), (252, 147, 7), (251, 146, 10), (252, 145, 7), (254, 148, 10), (254, 149, 25), (253, 148, 17), (254, 149, 13), (254, 152, 39), (252, 153, 42), (253, 153, 38), (253, 151, 38), (254, 151, 47), (253, 153, 46), (254, 154, 52), (254, 153, 46), (252, 154, 36), (254, 157, 52), (253, 159, 58), (253, 160, 62), (251, 160, 47), (254, 161, 59), (254, 161, 69), (253, 163, 69), (252, 166, 74), (252, 169, 78), (252, 172, 83), (253, 175, 87), (251, 176, 88), (253, 181, 107), (254, 183, 116), (253, 185, 115), (253, 185, 120), (253, 187, 126), (252, 190, 131), (252, 192, 138), (252, 192, 143), (252, 197, 151), (253, 207, 165), (252, 207, 168), (179, 44, 33), (169, 0, 0), (189, 25, 7), (182, 20, 1), (172, 5, 0), (169, 0, 2), (166, 0, 2), (162, 0, 1), (160, 0, 0), (159, 0, 1), (155, 1, 1), (154, 0, 1), (146, 2, 2), (189, 63, 21), (175, 7, 4), (177, 0, 1), (176, 0, 0), (178, 6, 3), (204, 35, 15), (219, 54, 25), (219, 57, 34), (221, 59, 40), (225, 64, 44), (224, 64, 38), (234, 21, 175), (238, 41, 130), (234, 66, 15), (239, 81, 12), (241, 90, 17), (240, 90, 29), (195, 18, 6), (195, 13, 0), (196, 22, 2), (189, 47, 6), (242, 189, 20), (232, 199, 7), (217, 177, 1), (211, 166, 1), (208, 159, 2), (209, 164, 1), (208, 172, 0), (198, 151, 28), (148, 46, 63), (122, 0, 40), (116, 0, 12), (131, 0, 0), (127, 6, 4), (111, 3, 12), (159, 12, 9), (239, 107, 40), (244, 128, 23), (219, 95, 1), (211, 85, 0), (207, 78, 1), (203, 72, 0), (200, 66, 0), (202, 66, 1), (202, 66, 2), (196, 63, 0), (214, 89, 4), (243, 127, 7), (239, 128, 7), (234, 120, 4), (236, 120, 2), (239, 120, 1), (243, 121, 1), (245, 123, 3), (246, 125, 3), (249, 127, 1), (252, 129, 2), (253, 131, 1), (253, 133, 1), (253, 135, 2), (254, 136, 2), (254, 139, 1), (255, 143, 2), (250, 130, 15), (158, 41, 6), (89, 17, 2), (97, 29, 20), (102, 31, 33), (96, 21, 37), (122, 64, 45), (230, 214, 99), (255, 255, 87), (255, 250, 56), (255, 247, 50), (255, 250, 72), (255, 255, 102), (224, 208, 110), (89, 60, 49), (111, 69, 60), (169, 133, 69), (239, 225, 97), (255, 249, 77), (255, 237, 43), (254, 233, 42), (255, 237, 62), (255, 244, 137), (255, 233, 216), (254, 218, 195), (254, 206, 162), (253, 198, 155), (253, 191, 146), (252, 187, 122), (251, 173, 101), (255, 170, 100), (253, 165, 85), (252, 160, 69), (253, 158, 66), (253, 155, 69), (253, 153, 65), (253, 150, 55), (252, 149, 40), (253, 144, 19), (253, 145, 15), (255, 147, 32), (254, 147, 39), (253, 147, 33), (254, 144, 17), (253, 141, 5), (252, 141, 3), (252, 140, 2), (253, 141, 2), (253, 143, 2), (254, 143, 2), (253, 142, 1), (255, 145, 2), (254, 148, 16), (253, 147, 25), (252, 147, 21), (253, 148, 18), (253, 147, 25), (252, 147, 21), (253, 148, 29), (253, 148, 27), (252, 149, 22), (255, 153, 45), (254, 153, 55), (255, 155, 55), (252, 154, 39), (255, 155, 50), (254, 157, 57), (253, 159, 59), (253, 162, 62), (253, 165, 69), (254, 166, 72), (253, 167, 71), (252, 167, 72), (254, 171, 101), (254, 174, 103), (253, 175, 101), (253, 178, 107), (253, 180, 113), (252, 183, 120), (254, 187, 124), (252, 187, 123), (250, 192, 137), (250, 197, 149), (254, 211, 162), (232, 159, 124), (167, 6, 4), (181, 13, 4), (175, 12, 4), (167, 1, 0), (162, 1, 1), (160, 0, 2), (158, 1, 1), (156, 0, 0), (155, 1, 2), (153, 1, 1), (147, 0, 2), (163, 31, 4), (239, 147, 19), (190, 42, 10), (169, 0, 0), (175, 0, 0), (199, 34, 12), (216, 66, 35), (215, 68, 43), (212, 66, 43), (209, 59, 34), (200, 41, 18), (197, 23, 0), (234, 0, 132), (232, 0, 124), (232, 32, 28), (224, 55, 0), (226, 59, 0), (225, 66, 4), (198, 29, 3), (193, 20, 5), (187, 46, 4), (217, 121, 14), (230, 180, 10), (220, 170, 2), (212, 162, 2), (202, 157, 2), (197, 152, 0), (201, 154, 2), (208, 168, 2), (171, 109, 21), (108, 0, 34), (126, 3, 21), (170, 31, 18), (194, 39, 9), (187, 28, 6), (154, 12, 8), (205, 84, 32), (241, 124, 21), (213, 87, 0), (209, 76, 4), (200, 65, 1), (195, 59, 2), (193, 55, 1), (191, 55, 1), (189, 53, 2), (188, 48, 3), (187, 52, 1), (226, 107, 8), (237, 123, 6), (233, 119, 5), (231, 114, 1), (232, 114, 1), (233, 114, 0), (235, 116, 0), (238, 117, 1), (241, 118, 2), (244, 120, 1), (247, 123, 2), (249, 125, 1), (250, 127, 1), (251, 129, 2), (253, 131, 2), (254, 134, 1), (253, 135, 1), (255, 144, 4), (220, 103, 11), (84, 9, 0), (83, 16, 9), (90, 19, 21), (99, 37, 20), (232, 198, 62), (255, 240, 27), (251, 220, 0), (255, 219, 0), (255, 219, 0), (253, 222, 0), (251, 225, 0), (255, 239, 40), (247, 238, 100), (255, 250, 139), (255, 247, 91), (255, 220, 20), (252, 210, 0), (252, 210, 0), (250, 211, 0), (247, 212, 3), (251, 222, 154), (253, 222, 211), (253, 208, 176), (255, 197, 152), (251, 190, 133), (252, 183, 125), (251, 174, 106), (250, 166, 85), (253, 162, 79), (253, 159, 73), (253, 157, 64), (253, 153, 61), (253, 150, 57), (254, 149, 52), (253, 146, 48), (253, 142, 24), (254, 142, 0), (253, 141, 11), (255, 142, 27), (254, 143, 17), (252, 141, 13), (254, 140, 18), (253, 138, 7), (253, 138, 1), (252, 137, 0), (253, 138, 0), (254, 140, 1), (254, 140, 0), (254, 138, 0), (255, 139, 1), (254, 143, 5), (253, 144, 9), (253, 144, 6), (253, 144, 3), (253, 143, 4), (252, 144, 3), (253, 145, 6), (254, 144, 15), (252, 145, 15), (254, 149, 25), (253, 151, 34), (254, 151, 41), (252, 147, 32), (255, 151, 50), (254, 153, 53), (254, 155, 55), (253, 157, 56), (253, 159, 66), (254, 162, 71), (253, 161, 62), (252, 162, 60), (254, 166, 83), (254, 170, 84), (253, 169, 85), (254, 173, 98), (253, 174, 97), (252, 178, 110), (252, 181, 114), (251, 180, 108), (251, 181, 117), (252, 187, 134), (252, 197, 146), (255, 211, 166), (200, 90, 62), (165, 0, 0), (169, 2, 4), (166, 1, 0), (159, 1, 1), (156, 1, 1), (154, 1, 0), (153, 0, 0), (154, 1, 2), (148, 0, 0), (148, 8, 10), (231, 156, 38), (244, 180, 3), (220, 110, 11), (190, 45, 31), (224, 95, 81), (245, 144, 120), (248, 159, 132), (251, 159, 132), (253, 158, 130), (249, 153, 121), (240, 136, 104), (225, 94, 73), (227, 28, 113), (225, 34, 102), (225, 50, 36), (219, 52, 2), (215, 38, 0), (211, 40, 0), (222, 74, 21), (246, 111, 43), (241, 129, 24), (230, 150, 4), (237, 146, 1), (248, 139, 2), (248, 137, 5), (226, 136, 6), (191, 137, 2), (184, 137, 2), (188, 143, 3), (160, 103, 10), (107, 3, 9), (173, 20, 10), (199, 29, 6), (191, 22, 0), (184, 11, 1), (200, 41, 9), (241, 114, 18), (214, 87, 0), (204, 71, 4), (197, 63, 3), (192, 56, 0), (189, 52, 0), (187, 51, 1), (184, 49, 1), (182, 46, 1), (179, 40, 1), (199, 69, 6), (232, 117, 7), (231, 117, 7), (226, 111, 3), (226, 108, 1), (226, 107, 0), (226, 107, 1), (227, 109, 1), (230, 110, 0), (233, 112, 0), (236, 114, 1), (239, 116, 1), (241, 118, 1), (242, 120, 0), (245, 119, 0), (246, 116, 0), (248, 117, 0), (249, 120, 0), (253, 125, 0), (238, 129, 8), (162, 115, 61), (193, 173, 106), (208, 193, 123), (216, 196, 87), (255, 221, 15), (254, 212, 0), (254, 210, 0), (253, 212, 0), (254, 212, 0), (255, 214, 0), (254, 216, 0), (252, 218, 0), (252, 232, 18), (255, 237, 33), (254, 213, 5), (255, 203, 0), (254, 199, 0), (254, 198, 0), (253, 196, 0), (251, 207, 77), (252, 217, 203), (249, 213, 181), (254, 198, 156), (255, 187, 135), (253, 179, 117), (252, 171, 103), (253, 165, 90), (252, 157, 71), (253, 154, 64), (253, 153, 61), (252, 149, 51), (251, 146, 43), (254, 146, 45), (255, 146, 47), (253, 144, 40), (253, 139, 19), (254, 138, 0), (253, 137, 8), (254, 138, 18), (252, 139, 4), (252, 138, 2), (253, 138, 5), (252, 135, 0), (253, 135, 0), (253, 136, 1), (253, 136, 1), (254, 136, 2), (254, 136, 1), (255, 136, 1), (254, 136, 2), (253, 139, 2), (253, 140, 1), (253, 140, 1), (253, 140, 2), (254, 141, 3), (254, 140, 3), (253, 140, 2), (254, 140, 6), (253, 142, 6), (252, 144, 5), (252, 146, 14), (253, 146, 17), (252, 144, 23), (255, 147, 47), (254, 150, 46), (254, 152, 51), (252, 153, 49), (253, 155, 60), (255, 158, 68), (253, 157, 50), (253, 159, 51), (254, 162, 68), (255, 164, 68), (253, 164, 68), (254, 167, 74), (251, 167, 74), (252, 170, 89), (253, 177, 105), (252, 175, 101), (252, 174, 101), (252, 180, 121), (251, 190, 140), (252, 200, 152), (250, 191, 124), (205, 108, 23), (163, 25, 4), (150, 0, 2), (155, 0, 3), (155, 0, 0), (150, 0, 1), (146, 0, 0), (141, 0, 0), (150, 13, 5), (220, 132, 27), (252, 213, 16), (241, 176, 27), (246, 155, 86), (255, 158, 140), (255, 154, 133), (252, 141, 117), (251, 128, 105), (251, 122, 99), (254, 120, 99), (254, 121, 97), (255, 129, 104), (255, 140, 115), (251, 171, 84), (253, 174, 81), (250, 171, 68), (243, 154, 62), (232, 115, 40), (208, 57, 8), (228, 77, 6), (255, 124, 13), (252, 115, 10), (252, 120, 5), (251, 116, 2), (250, 110, 1), (247, 106, 0), (243, 106, 3), (219, 115, 3), (176, 128, 0), (171, 130, 0), (175, 124, 14), (180, 81, 69), (176, 17, 17), (169, 0, 0), (163, 0, 0), (157, 0, 2), (203, 59, 10), (227, 97, 4), (207, 72, 2), (199, 61, 4), (191, 54, 0), (189, 51, 0), (187, 48, 0), (185, 48, 0), (183, 47, 0), (181, 45, 1), (177, 39, 2), (209, 84, 9), (232, 118, 8), (228, 113, 7), (220, 105, 2), (222, 102, 1), (223, 102, 0), (222, 103, 0), (222, 103, 0), (224, 104, 0), (226, 106, 0), (230, 108, 1), (234, 110, 1), (234, 111, 0), (234, 104, 0), (230, 126, 19), (237, 172, 66), (244, 192, 87), (244, 178, 79), (234, 146, 36), (240, 192, 62), (255, 251, 105), (255, 255, 79), (255, 254, 87), (255, 240, 57), (254, 208, 3), (254, 206, 0), (253, 206, 0), (254, 207, 0), (254, 209, 0), (254, 211, 0), (253, 211, 1), (253, 214, 1), (255, 216, 2), (254, 214, 0), (254, 205, 0), (255, 198, 0), (253, 195, 0), (253, 192, 0), (251, 195, 16), (254, 210, 154), (252, 209, 182), (251, 203, 165), (253, 190, 147), (254, 178, 121), (251, 170, 106), (251, 164, 90), (252, 158, 76), (251, 150, 50), (253, 148, 54), (254, 146, 58), (254, 144, 51), (252, 142, 29), (253, 142, 26), (253, 142, 27), (251, 141, 10), (253, 139, 4), (254, 135, 1), (253, 135, 1), (253, 135, 3), (252, 135, 1), (252, 135, 2), (253, 134, 1), (252, 132, 0), (253, 132, 1), (253, 132, 1), (254, 133, 1), (254, 133, 1), (253, 132, 0), (254, 133, 1), (253, 134, 2), (252, 136, 2), (252, 136, 0), (252, 136, 0), (252, 136, 0), (254, 137, 2), (255, 137, 2), (254, 137, 1), (253, 137, 1), (253, 139, 2), (253, 141, 1), (253, 142, 3), (252, 142, 1), (253, 143, 11), (255, 145, 29), (255, 147, 39), (254, 148, 46), (253, 149, 42), (254, 151, 53), (255, 152, 61), (251, 152, 43), (254, 155, 52), (254, 158, 63), (255, 158, 62), (253, 158, 58), (254, 161, 64), (252, 162, 67), (252, 163, 72), (252, 171, 93), (252, 173, 96), (250, 171, 88), (251, 176, 109), (252, 180, 122), (254, 188, 135), (255, 198, 153), (231, 180, 70), (209, 126, 6), (175, 49, 13), (149, 8, 7), (142, 0, 3), (140, 0, 3), (147, 11, 6), (173, 56, 10), (225, 139, 11), (243, 186, 3), (242, 167, 37), (254, 144, 113), (255, 131, 116), (254, 114, 90), (251, 100, 72), (251, 93, 64), (250, 91, 57), (250, 89, 55), (251, 88, 56), (251, 90, 59), (252, 89, 60), (253, 95, 66), (254, 156, 4), (254, 156, 4), (252, 159, 8), (252, 164, 22), (255, 173, 38), (250, 158, 37), (243, 129, 18), (243, 101, 2), (242, 98, 0), (243, 98, 4), (239, 92, 4), (233, 87, 3), (228, 82, 1), (222, 77, 2), (217, 81, 4), (200, 133, 4), (178, 134, 4), (188, 127, 79), (195, 91, 110), (166, 9, 12), (169, 5, 5), (169, 11, 9), (157, 4, 3), (203, 65, 9), (215, 81, 1), (202, 63, 1), (196, 54, 1), (190, 48, 0), (189, 47, 0), (186, 46, 0), (183, 45, 1), (181, 45, 1), (178, 44, 2), (176, 41, 4), (213, 92, 9), (228, 116, 9), (220, 104, 2), (216, 99, 1), (217, 99, 0), (218, 98, 0), (217, 99, 0), (219, 98, 0), (219, 99, 0), (220, 100, 0), (222, 102, 0), (225, 103, 0), (225, 96, 0), (230, 146, 43), (248, 228, 124), (252, 246, 130), (249, 250, 121), (247, 252, 123), (247, 248, 127), (252, 249, 148), (251, 247, 142), (249, 241, 91), (246, 232, 29), (252, 216, 0), (254, 202, 0), (250, 204, 6), (249, 211, 17), (251, 211, 16), (249, 208, 7), (252, 204, 0), (254, 205, 0), (253, 207, 0), (255, 209, 2), (253, 203, 1), (252, 197, 0), (253, 196, 0), (254, 194, 1), (250, 192, 0), (247, 203, 74), (254, 207, 176), (253, 196, 155), (253, 190, 141), (254, 179, 125), (254, 167, 103), (251, 162, 86), (252, 156, 69), (253, 150, 64), (250, 144, 35), (253, 147, 43), (254, 143, 38), (255, 141, 37), (253, 138, 27), (254, 138, 22), (254, 138, 19), (253, 136, 5), (254, 135, 2), (253, 132, 1), (252, 131, 0), (253, 132, 0), (253, 132, 0), (253, 132, 1), (253, 132, 1), (253, 131, 1), (253, 129, 0), (254, 129, 0), (254, 130, 0), (254, 131, 0), (254, 130, 0), (253, 131, 0), (253, 132, 0), (252, 133, 1), (253, 133, 0), (253, 133, 0), (253, 133, 0), (253, 133, 0), (254, 134, 1), (254, 132, 0), (254, 135, 1), (254, 138, 2), (253, 137, 2), (253, 137, 0), (253, 137, 2), (253, 140, 5), (253, 143, 5), (253, 144, 12), (252, 145, 20), (254, 148, 25), (255, 148, 35), (254, 149, 41), (249, 147, 31), (253, 151, 47), (254, 153, 54), (254, 155, 54), (254, 155, 52), (253, 155, 54), (251, 155, 52), (254, 160, 66), (251, 165, 83), (252, 167, 88), (252, 167, 85), (253, 169, 92), (251, 170, 99), (251, 179, 115), (253, 192, 146), (242, 189, 126), (212, 145, 13), (221, 148, 8), (207, 129, 12), (195, 113, 12), (200, 116, 14), (216, 126, 15), (226, 147, 8), (230, 155, 0), (237, 148, 24), (253, 132, 106), (254, 111, 93), (251, 91, 63), (253, 78, 43), (250, 72, 29), (249, 66, 21), (248, 64, 15), (249, 63, 13), (249, 63, 16), (247, 67, 20), (248, 68, 24), (251, 74, 36), (253, 131, 0), (254, 130, 0), (253, 129, 1), (253, 130, 0), (253, 135, 0), (251, 147, 6), (254, 155, 15), (251, 139, 22), (238, 99, 7), (227, 79, 0), (226, 73, 0), (223, 67, 0), (218, 63, 0), (211, 59, 1), (201, 60, 1), (209, 132, 3), (202, 143, 48), (176, 88, 103), (176, 62, 78), (203, 51, 20), (217, 55, 12), (217, 59, 12), (210, 47, 7), (211, 65, 5), (205, 69, 4), (198, 56, 4), (193, 49, 0), (189, 44, 0), (188, 44, 1), (182, 44, 0), (180, 45, 1), (178, 46, 2), (175, 44, 1), (173, 44, 0), (217, 98, 11), (225, 111, 8), (214, 100, 0), (213, 91, 0), (212, 82, 0), (211, 83, 0), (207, 85, 0), (211, 85, 0), (212, 85, 0), (212, 87, 0), (214, 93, 0), (218, 91, 0), (219, 125, 18), (249, 229, 67), (253, 230, 34), (252, 220, 7), (251, 221, 4), (253, 224, 7), (255, 228, 17), (251, 237, 61), (250, 248, 132), (252, 248, 167), (252, 247, 142), (246, 226, 61), (250, 222, 74), (251, 239, 127), (250, 247, 150), (253, 247, 147), (250, 242, 125), (246, 226, 76), (250, 205, 13), (255, 203, 0), (255, 205, 2), (254, 200, 1), (254, 195, 0), (254, 194, 0), (255, 193, 0), (253, 194, 12), (253, 200, 132), (254, 197, 160), (254, 188, 143), (253, 177, 119), (253, 169, 97), (254, 160, 79), (254, 154, 67), (253, 148, 53), (253, 146, 54), (252, 142, 36), (255, 144, 38), (253, 138, 14), (254, 136, 11), (253, 136, 16), (253, 135, 12), (253, 135, 6), (254, 135, 2), (254, 132, 1), (253, 130, 1), (252, 129, 0), (254, 130, 0), (254, 130, 0), (254, 130, 1), (255, 130, 2), (255, 129, 2), (255, 128, 0), (255, 128, 0), (254, 129, 1), (254, 129, 1), (253, 129, 0), (254, 129, 1), (254, 130, 1), (254, 131, 1), (254, 132, 0), (254, 132, 0), (254, 132, 0), (254, 132, 0), (253, 131, 0), (254, 130, 1), (254, 131, 1), (254, 134, 2), (254, 134, 2), (253, 134, 1), (253, 135, 2), (253, 137, 2), (253, 139, 0), (252, 140, 0), (252, 141, 3), (254, 143, 14), (255, 144, 20), (254, 145, 23), (252, 144, 29), (253, 145, 36), (254, 147, 38), (253, 150, 41), (254, 151, 53), (254, 153, 50), (252, 151, 39), (254, 155, 54), (251, 159, 67), (252, 162, 74), (251, 164, 82), (253, 167, 87), (253, 169, 95), (251, 173, 108), (249, 180, 119), (254, 195, 146), (219, 153, 45), (209, 141, 0), (216, 151, 1), (218, 158, 4), (217, 154, 2), (215, 133, 1), (214, 133, 0), (219, 127, 17), (250, 124, 87), (254, 103, 74), (248, 83, 40), (243, 68, 24), (245, 57, 7), (241, 53, 1), (241, 50, 0), (242, 47, 0), (243, 45, 0), (242, 46, 0), (240, 49, 0), (241, 52, 5), (245, 57, 9), (249, 120, 0), (253, 118, 2), (253, 117, 1), (251, 118, 0), (251, 120, 0), (253, 121, 0), (254, 124, 0), (255, 139, 9), (251, 123, 15), (231, 83, 1), (229, 77, 1), (229, 75, 3), (222, 72, 3), (205, 59, 1), (188, 63, 0), (185, 122, 4), (176, 111, 65), (162, 60, 81), (194, 52, 34), (209, 48, 5), (203, 40, 0), (197, 37, 0), (196, 33, 0), (205, 55, 3), (200, 59, 1), (194, 50, 3), (190, 44, 1), (188, 41, 0), (185, 40, 0), (180, 41, 0), (178, 44, 2), (178, 45, 4), (175, 44, 3), (170, 41, 5), (217, 96, 13), (215, 96, 0), (211, 92, 0), (210, 117, 25), (220, 146, 69), (226, 170, 95), (228, 179, 110), (231, 178, 107), (225, 167, 94), (223, 140, 69), (214, 112, 24), (210, 81, 0), (234, 162, 17), (255, 223, 10), (253, 210, 0), (252, 211, 0), (252, 211, 0), (250, 213, 0), (249, 226, 22), (249, 243, 114), (250, 248, 167), (252, 245, 167), (254, 248, 157), (254, 245, 140), (253, 240, 109), (254, 240, 87), (252, 239, 75), (253, 239, 77), (252, 244, 96), (253, 248, 123), (253, 234, 105), (246, 209, 22), (253, 201, 1), (253, 201, 3), (250, 201, 11), (251, 201, 18), (248, 200, 3), (249, 198, 56), (254, 195, 151), (251, 191, 138), (252, 182, 128), (255, 169, 106), (253, 164, 88), (253, 155, 72), (254, 148, 57), (252, 144, 51), (250, 144, 48), (251, 139, 27), (252, 134, 16), (250, 132, 8), (251, 131, 2), (252, 132, 5), (252, 131, 3), (254, 131, 1), (253, 131, 1), (253, 129, 0), (253, 127, 0), (253, 127, 0), (255, 127, 0), (254, 126, 0), (253, 126, 0), (253, 125, 1), (253, 125, 1), (253, 125, 1), (253, 125, 1), (253, 125, 1), (254, 126, 1), (254, 125, 0), (255, 126, 2), (254, 128, 1), (254, 128, 0), (254, 128, 0), (254, 128, 0), (254, 128, 0), (254, 128, 1), (254, 128, 1), (254, 128, 0), (254, 128, 1), (254, 129, 2), (254, 130, 2), (252, 131, 1), (254, 133, 1), (254, 134, 1), (254, 135, 0), (254, 137, 2), (254, 138, 1), (254, 138, 4), (255, 139, 7), (253, 140, 7), (251, 141, 11), (252, 141, 23), (253, 143, 25), (254, 145, 35), (254, 147, 49), (252, 149, 39), (252, 149, 32), (254, 152, 50), (252, 154, 63), (252, 157, 68), (251, 161, 79), (251, 163, 81), (253, 167, 90), (255, 170, 103), (249, 174, 109), (254, 193, 146), (238, 174, 86), (204, 139, 1), (208, 145, 1), (207, 147, 2), (207, 143, 3), (205, 125, 3), (205, 119, 2), (229, 117, 49), (254, 98, 75), (248, 71, 29), (245, 58, 12), (238, 49, 4), (237, 43, 0), (237, 39, 0), (236, 36, 0), (236, 34, 0), (236, 34, 0), (236, 34, 1), (237, 37, 1), (237, 38, 1), (238, 42, 1), (245, 109, 3), (246, 109, 3), (244, 107, 1), (244, 108, 1), (246, 107, 1), (247, 107, 1), (248, 106, 0), (249, 112, 0), (254, 122, 6), (241, 100, 4), (229, 83, 2), (233, 91, 4), (243, 108, 14), (224, 88, 13), (187, 59, 1), (185, 77, 5), (170, 62, 43), (168, 44, 43), (194, 26, 5), (186, 17, 0), (177, 10, 0), (170, 8, 0), (163, 1, 0), (179, 25, 3), (198, 53, 3), (190, 44, 1), (187, 39, 0), (184, 37, 0), (181, 38, 0), (179, 38, 0), (179, 41, 3), (177, 42, 4), (174, 40, 3), (172, 35, 1), (203, 82, 12), (221, 147, 59), (235, 206, 140), (248, 243, 201), (255, 255, 220), (255, 255, 225), (255, 255, 225), (255, 255, 219), (255, 255, 218), (254, 255, 214), (249, 242, 186), (234, 197, 132), (242, 203, 57), (250, 210, 0), (253, 206, 0), (254, 207, 1), (252, 204, 0), (248, 216, 31), (253, 240, 146), (254, 239, 172), (252, 236, 145), (253, 236, 141), (252, 236, 113), (250, 227, 47), (252, 219, 6), (252, 220, 0), (252, 220, 0), (252, 221, 0), (252, 224, 3), (252, 228, 14), (249, 239, 65), (250, 229, 71), (246, 205, 5), (252, 218, 25), (254, 230, 64), (254, 234, 78), (252, 232, 62), (250, 206, 128), (252, 187, 141), (253, 181, 120), (249, 171, 110), (254, 161, 93), (253, 155, 76), (252, 150, 62), (254, 145, 56), (254, 142, 51), (249, 139, 36), (251, 134, 13), (253, 131, 2), (252, 131, 4), (253, 129, 3), (253, 129, 2), (253, 128, 0), (254, 128, 0), (254, 127, 0), (253, 125, 0), (252, 123, 0), (253, 123, 0), (254, 124, 0), (253, 123, 0), (252, 122, 0), (252, 121, 0), (252, 121, 0), (253, 122, 1), (253, 122, 1), (253, 122, 1), (254, 123, 0), (255, 123, 0), (255, 124, 1), (255, 126, 0), (254, 126, 0), (254, 125, 1), (254, 125, 1), (254, 125, 1), (253, 125, 1), (253, 125, 1), (254, 125, 1), (254, 126, 1), (255, 126, 1), (253, 128, 0), (251, 128, 0), (253, 131, 1), (254, 131, 1), (254, 132, 1), (255, 133, 3), (255, 135, 2), (255, 135, 0), (254, 136, 0), (254, 136, 0), (253, 137, 0), (253, 139, 6), (253, 140, 18), (255, 142, 34), (253, 144, 36), (250, 145, 21), (253, 146, 30), (254, 150, 46), (254, 151, 52), (253, 154, 65), (253, 159, 70), (251, 158, 70), (253, 163, 80), (254, 166, 90), (250, 170, 102), (253, 183, 133), (248, 182, 121), (203, 145, 16), (201, 143, 0), (203, 146, 2), (207, 146, 7), (201, 123, 1), (210, 114, 13), (242, 104, 55), (247, 72, 25), (243, 51, 6), (240, 40, 1), (236, 35, 1), (234, 30, 2), (233, 27, 5), (234, 24, 4), (233, 22, 4), (234, 23, 4), (233, 24, 5), (234, 26, 5), (234, 30, 2), (232, 33, 1), (237, 103, 2), (237, 101, 2), (237, 101, 2), (236, 100, 1), (236, 99, 0), (236, 99, 0), (237, 97, 1), (239, 98, 2), (245, 107, 1), (236, 92, 6), (209, 56, 2), (209, 60, 2), (201, 54, 6), (191, 32, 3), (194, 25, 2), (196, 20, 2), (189, 13, 0), (179, 7, 0), (175, 0, 0), (172, 0, 2), (169, 0, 2), (163, 0, 0), (155, 0, 0), (154, 3, 1), (186, 36, 8), (190, 42, 4), (183, 36, 0), (182, 36, 1), (180, 36, 2), (177, 35, 0), (177, 38, 2), (177, 39, 3), (169, 22, 0), (184, 77, 33), (227, 199, 143), (255, 255, 206), (252, 255, 206), (253, 247, 192), (250, 244, 184), (250, 244, 180), (252, 243, 176), (253, 244, 175), (251, 246, 177), (252, 247, 177), (253, 251, 190), (254, 255, 211), (254, 255, 204), (249, 234, 122), (246, 210, 18), (252, 202, 0), (251, 206, 6), (251, 225, 73), (253, 218, 82), (254, 206, 50), (253, 207, 37), (252, 218, 45), (250, 218, 26), (252, 208, 0), (253, 206, 0), (252, 205, 0), (255, 204, 0), (252, 208, 0), (254, 209, 0), (255, 211, 0), (252, 218, 2), (254, 224, 39), (252, 221, 19), (254, 220, 7), (254, 221, 17), (252, 223, 17), (252, 220, 49), (248, 198, 138), (249, 180, 120), (252, 172, 111), (249, 167, 101), (251, 156, 82), (251, 149, 65), (253, 144, 56), (250, 141, 51), (251, 137, 31), (251, 132, 21), (252, 131, 12), (253, 129, 3), (253, 128, 4), (253, 126, 2), (254, 125, 1), (253, 124, 0), (253, 124, 0), (254, 123, 0), (253, 123, 1), (253, 121, 0), (254, 121, 0), (254, 121, 1), (253, 121, 0), (254, 119, 0), (254, 118, 0), (252, 119, 0), (254, 120, 0), (254, 120, 1), (254, 120, 2), (255, 122, 1), (254, 122, 1), (255, 122, 1), (255, 123, 1), (254, 123, 1), (254, 122, 1), (254, 122, 1), (254, 122, 1), (254, 122, 1), (254, 122, 1), (255, 123, 1), (254, 123, 1), (253, 125, 1), (254, 127, 2), (253, 126, 1), (255, 127, 2), (254, 128, 1), (255, 129, 1), (255, 130, 1), (255, 131, 1), (254, 131, 0), (254, 132, 0), (254, 133, 0), (254, 134, 2), (253, 136, 3), (253, 137, 10), (254, 138, 22), (254, 140, 24), (251, 141, 14), (252, 142, 19), (253, 145, 26), (252, 147, 30), (252, 150, 48), (253, 153, 61), (252, 154, 65), (254, 159, 75), (253, 160, 79), (253, 166, 97), (251, 174, 120), (254, 182, 129), (216, 154, 36), (199, 141, 0), (203, 146, 5), (202, 136, 5), (201, 117, 0), (221, 114, 20), (244, 77, 35), (240, 51, 6), (234, 40, 4), (230, 29, 2), (229, 23, 2), (225, 13, 0), (228, 7, 1), (231, 6, 1), (232, 4, 0), (232, 4, 0), (231, 5, 1), (231, 10, 2), (231, 16, 1), (229, 24, 0), (230, 95, 0), (230, 95, 0), (231, 95, 0), (231, 95, 0), (232, 93, 0), (231, 91, 0), (231, 89, 0), (232, 89, 0), (237, 92, 1), (236, 89, 10), (204, 49, 6), (198, 38, 9), (176, 6, 0), (177, 0, 1), (179, 0, 1), (173, 0, 0), (175, 0, 0), (175, 5, 4), (174, 8, 6), (167, 3, 3), (159, 0, 0), (154, 0, 2), (148, 0, 0), (142, 0, 0), (158, 7, 2), (183, 35, 5), (183, 34, 0), (180, 32, 1), (179, 32, 1), (175, 33, 0), (176, 35, 1), (166, 25, 0), (183, 89, 44), (246, 230, 172), (255, 255, 198), (252, 238, 168), (253, 235, 156), (253, 235, 148), (252, 234, 141), (253, 233, 137), (254, 233, 137), (254, 233, 138), (254, 234, 140), (254, 236, 142), (255, 239, 154), (255, 242, 168), (254, 245, 185), (253, 253, 199), (249, 246, 160), (248, 211, 31), (253, 199, 4), (253, 210, 19), (250, 193, 3), (253, 185, 0), (252, 183, 0), (253, 204, 6), (255, 203, 3), (255, 196, 1), (254, 194, 0), (253, 191, 0), (254, 190, 0), (255, 196, 2), (254, 200, 1), (253, 203, 1), (254, 207, 0), (255, 212, 5), (254, 213, 10), (251, 207, 0), (251, 203, 0), (250, 203, 0), (251, 201, 52), (251, 188, 136), (251, 170, 104), (254, 164, 93), (253, 159, 88), (252, 149, 73), (253, 143, 56), (252, 138, 32), (251, 134, 20), (252, 129, 17), (252, 129, 15), (252, 128, 12), (249, 125, 3), (251, 123, 2), (252, 122, 2), (253, 123, 1), (252, 121, 0), (252, 121, 1), (252, 120, 1), (253, 121, 1), (254, 119, 0), (253, 119, 0), (252, 119, 1), (253, 119, 0), (252, 117, 0), (252, 117, 0), (251, 118, 0), (253, 119, 1), (253, 119, 1), (254, 119, 2), (255, 120, 1), (253, 120, 1), (253, 120, 1), (254, 121, 1), (255, 122, 1), (255, 122, 1), (255, 122, 1), (255, 122, 1), (255, 121, 1), (255, 122, 1), (254, 121, 0), (252, 121, 0), (252, 122, 0), (254, 124, 2), (254, 124, 1), (254, 124, 1), (255, 126, 0), (255, 128, 0), (255, 128, 0), (255, 128, 0), (254, 128, 0), (253, 129, 0), (253, 130, 1), (254, 132, 2), (253, 132, 2), (254, 133, 3), (254, 136, 5), (252, 136, 6), (253, 138, 13), (252, 140, 7), (252, 140, 9), (254, 142, 30), (254, 146, 37), (252, 150, 48), (252, 151, 53), (254, 154, 70), (255, 157, 77), (253, 161, 90), (250, 165, 102), (255, 178, 119), (227, 161, 60), (196, 140, 0), (200, 143, 4), (196, 123, 1), (203, 122, 2), (223, 109, 16), (238, 59, 19), (232, 39, 2), (231, 26, 3), (230, 14, 1), (225, 5, 0), (224, 2, 1), (226, 0, 1), (227, 0, 0), (228, 0, 0), (228, 0, 0), (228, 0, 0), (227, 1, 0), (227, 1, 0), (230, 8, 1), (224, 88, 0), (224, 88, 1), (227, 89, 0), (228, 91, 0), (229, 90, 1), (228, 85, 1), (227, 82, 1), (228, 81, 0), (232, 80, 1), (234, 85, 3), (214, 67, 3), (184, 23, 4), (164, 0, 0), (167, 0, 0), (186, 32, 20), (211, 83, 44), (234, 116, 61), (240, 124, 64), (242, 121, 59), (234, 107, 46), (216, 86, 37), (203, 68, 37), (187, 49, 37), (170, 34, 30), (150, 17, 16), (153, 16, 7), (174, 28, 6), (177, 29, 5), (177, 28, 1), (174, 32, 0), (168, 21, 0), (180, 77, 34), (246, 235, 164), (255, 244, 171), (253, 230, 145), (249, 227, 123), (253, 223, 117), (255, 222, 108), (255, 221, 102), (255, 220, 99), (253, 222, 98), (255, 224, 101), (255, 225, 104), (254, 227, 106), (255, 229, 118), (254, 232, 131), (254, 237, 142), (255, 242, 155), (255, 248, 187), (253, 242, 154), (248, 205, 28), (253, 196, 0), (253, 186, 0), (252, 180, 0), (252, 177, 0), (253, 194, 3), (255, 198, 4), (255, 192, 1), (255, 190, 0), (255, 187, 0), (253, 187, 1), (254, 190, 2), (254, 193, 3), (253, 196, 2), (252, 199, 0), (254, 204, 2), (254, 201, 3), (252, 191, 0), (253, 188, 0), (252, 188, 0), (254, 186, 81), (253, 176, 124), (253, 162, 86), (255, 154, 77), (255, 151, 73), (254, 144, 60), (253, 137, 46), (252, 134, 21), (252, 131, 11), (252, 128, 18), (250, 126, 8), (251, 125, 8), (250, 121, 2), (249, 120, 1), (251, 120, 1), (251, 119, 0), (251, 119, 0), (250, 119, 1), (251, 118, 1), (252, 118, 0), (253, 117, 0), (251, 116, 0), (250, 117, 0), (250, 117, 0), (249, 116, 0), (249, 115, 0), (249, 115, 0), (252, 117, 2), (253, 117, 2), (253, 117, 1), (253, 117, 0), (253, 118, 0), (252, 118, 1), (252, 118, 0), (254, 120, 1), (254, 121, 0), (254, 121, 0), (254, 120, 2), (253, 119, 1), (253, 119, 0), (254, 121, 0), (254, 121, 0), (253, 121, 0), (254, 122, 1), (254, 122, 1), (254, 122, 0), (254, 123, 0), (253, 125, 0), (254, 125, 0), (254, 125, 0), (254, 125, 0), (253, 126, 1), (252, 128, 0), (254, 129, 1), (253, 129, 1), (254, 130, 0), (254, 132, 0), (253, 133, 3), (254, 136, 9), (255, 137, 8), (252, 137, 4), (253, 140, 12), (254, 143, 16), (254, 145, 26), (253, 146, 38), (254, 149, 60), (253, 153, 64), (253, 156, 74), (251, 157, 78), (255, 165, 95), (238, 166, 87), (194, 145, 3), (198, 136, 4), (197, 116, 2), (204, 130, 6), (218, 103, 5), (229, 48, 9), (229, 31, 4), (228, 11, 1), (226, 0, 0), (225, 0, 1), (227, 1, 2), (225, 2, 1), (226, 0, 0), (226, 0, 0), (226, 1, 0), (228, 1, 0), (228, 1, 0), (228, 1, 0), (229, 2, 2), (221, 84, 1), (221, 84, 2), (223, 87, 1), (225, 88, 0), (224, 84, 0), (224, 80, 0), (224, 76, 0), (225, 75, 0), (226, 72, 0), (233, 83, 1), (255, 122, 14), (239, 101, 13), (203, 55, 12), (219, 89, 52), (254, 148, 78), (255, 152, 62), (255, 140, 42), (249, 129, 24), (249, 124, 17), (249, 120, 15), (249, 119, 18), (247, 116, 20), (235, 100, 29), (203, 71, 38), (179, 46, 36), (165, 29, 25), (159, 18, 10), (166, 20, 5), (174, 27, 5), (175, 26, 0), (170, 43, 10), (240, 202, 137), (255, 240, 159), (254, 219, 125), (252, 215, 99), (252, 215, 87), (252, 213, 82), (254, 212, 74), (255, 210, 70), (255, 210, 68), (253, 212, 65), (253, 215, 68), (252, 217, 71), (252, 219, 76), (252, 221, 84), (251, 225, 93), (252, 229, 102), (253, 232, 122), (252, 237, 140), (251, 244, 161), (251, 217, 83), (249, 186, 1), (254, 179, 0), (253, 177, 0), (253, 174, 0), (253, 187, 2), (254, 195, 3), (254, 192, 0), (254, 190, 0), (254, 188, 3), (253, 188, 3), (253, 188, 1), (254, 190, 3), (254, 192, 3), (252, 195, 0), (253, 198, 2), (253, 190, 2), (253, 180, 0), (254, 179, 0), (251, 179, 12), (254, 180, 101), (255, 161, 103), (254, 153, 72), (253, 147, 68), (254, 145, 65), (253, 142, 54), (251, 136, 44), (252, 133, 29), (250, 128, 12), (250, 124, 8), (249, 122, 4), (250, 121, 3), (251, 120, 2), (250, 119, 2), (250, 118, 1), (250, 116, 0), (250, 116, 0), (251, 117, 1), (251, 118, 1), (250, 116, 0), (250, 116, 0), (250, 116, 0), (249, 115, 0), (249, 115, 0), (250, 115, 0), (251, 114, 2), (251, 114, 2), (252, 115, 2), (252, 115, 2), (251, 115, 1), (251, 114, 0), (251, 114, 0), (252, 116, 0), (253, 117, 1), (254, 118, 1), (254, 118, 1), (254, 118, 1), (254, 118, 1), (254, 118, 2), (254, 118, 1), (254, 118, 0), (254, 118, 0), (254, 118, 1), (255, 119, 2), (255, 119, 1), (253, 121, 1), (253, 122, 1), (254, 121, 1), (255, 121, 0), (255, 122, 0), (255, 123, 1), (255, 124, 2), (253, 126, 0), (254, 128, 1), (254, 128, 1), (254, 128, 1), (254, 128, 1), (253, 128, 1), (254, 130, 3), (255, 133, 5), (254, 135, 4), (254, 136, 4), (255, 139, 7), (253, 142, 11), (254, 143, 30), (254, 146, 46), (253, 148, 54), (253, 151, 67), (252, 153, 66), (255, 158, 80), (240, 160, 101), (103, 71, 18), (134, 82, 11), (207, 126, 6), (206, 132, 7), (215, 105, 4), (224, 39, 2), (227, 22, 1), (226, 3, 1), (225, 0, 1), (225, 0, 1), (226, 0, 1), (226, 0, 1), (226, 0, 1), (226, 0, 1), (226, 0, 1), (226, 0, 1), (226, 0, 1), (227, 1, 2), (227, 1, 2), (216, 80, 0), (219, 82, 1), (221, 84, 1), (218, 81, 0), (219, 78, 0), (220, 77, 0), (222, 75, 0), (223, 74, 1), (222, 72, 0), (232, 82, 3), (252, 109, 6), (251, 127, 11), (255, 149, 49), (255, 146, 56), (249, 131, 35), (243, 117, 14), (244, 108, 3), (243, 104, 0), (239, 101, 0), (236, 97, 0), (235, 96, 0), (234, 96, 0), (237, 100, 0), (231, 96, 12), (186, 54, 13), (146, 14, 8), (139, 7, 4), (138, 3, 1), (143, 6, 3), (140, 5, 0), (204, 129, 71), (255, 238, 153), (255, 211, 112), (253, 206, 84), (252, 201, 63), (253, 199, 56), (255, 198, 52), (255, 199, 42), (254, 200, 29), (254, 201, 29), (254, 201, 27), (254, 202, 29), (254, 204, 35), (254, 208, 40), (254, 210, 48), (254, 212, 57), (255, 217, 65), (255, 220, 86), (254, 224, 104), (253, 229, 111), (253, 217, 75), (251, 175, 6), (253, 171, 3), (254, 175, 2), (253, 175, 1), (252, 178, 1), (253, 193, 3), (252, 195, 1), (253, 192, 0), (253, 189, 2), (254, 189, 2), (253, 189, 1), (254, 191, 2), (254, 192, 1), (252, 195, 0), (254, 194, 3), (254, 178, 2), (254, 173, 0), (254, 173, 0), (250, 176, 26), (254, 172, 105), (254, 154, 84), (253, 147, 60), (251, 143, 56), (252, 140, 53), (252, 139, 49), (251, 135, 40), (251, 130, 26), (251, 126, 13), (249, 123, 3), (250, 120, 2), (251, 119, 1), (250, 119, 0), (249, 117, 0), (250, 115, 0), (249, 116, 0), (249, 116, 1), (250, 116, 1), (250, 116, 0), (249, 115, 0), (249, 115, 0), (249, 115, 0), (248, 113, 0), (249, 112, 0), (249, 113, 2), (249, 113, 3), (250, 113, 2), (250, 114, 1), (250, 114, 1), (250, 114, 1), (249, 113, 1), (249, 113, 0), (251, 115, 0), (252, 116, 0), (253, 117, 1), (253, 117, 2), (253, 117, 2), (253, 117, 1), (252, 116, 0), (252, 116, 0), (253, 117, 0), (253, 117, 1), (253, 117, 2), (253, 116, 2), (253, 117, 0), (252, 118, 0), (252, 119, 1), (253, 119, 1), (253, 118, 1), (252, 119, 0), (254, 121, 0), (254, 121, 0), (253, 122, 0), (253, 125, 0), (254, 125, 1), (254, 125, 1), (253, 124, 0), (253, 125, 0), (255, 127, 1), (255, 130, 2), (254, 132, 2), (255, 134, 3), (254, 135, 3), (252, 137, 3), (253, 139, 15), (252, 142, 36), (252, 143, 45), (254, 147, 61), (253, 148, 66), (253, 150, 70), (247, 152, 80), (73, 41, 29), (109, 68, 9), (213, 132, 4), (204, 131, 5), (210, 119, 5), (220, 40, 6), (228, 11, 1), (226, 1, 0), (225, 1, 1), (225, 0, 1), (226, 0, 1), (226, 0, 1), (227, 1, 2), (227, 1, 2), (226, 0, 1), (226, 0, 1), (226, 0, 1), (226, 0, 1), (226, 0, 1), (215, 79, 0), (219, 81, 2), (217, 78, 1), (214, 75, 1), (217, 75, 1), (219, 75, 1), (223, 74, 2), (224, 73, 3), (223, 70, 2), (227, 68, 0), (236, 81, 5), (250, 125, 45), (248, 133, 39), (242, 115, 9), (237, 105, 1), (237, 102, 0), (237, 98, 0), (238, 96, 0), (236, 94, 0), (233, 92, 0), (232, 91, 1), (228, 88, 3), (226, 86, 4), (227, 89, 0), (218, 87, 6), (153, 22, 2), (123, 0, 0), (128, 2, 2), (124, 0, 1), (125, 14, 13), (239, 198, 117), (255, 217, 112), (253, 201, 78), (253, 195, 49), (253, 192, 32), (255, 189, 26), (255, 186, 20), (254, 188, 11), (254, 191, 4), (254, 191, 4), (255, 191, 4), (254, 192, 3), (253, 194, 4), (253, 198, 8), (254, 200, 13), (252, 203, 20), (253, 208, 28), (254, 211, 51), (255, 212, 63), (250, 214, 62), (253, 210, 41), (252, 176, 2), (250, 161, 3), (252, 169, 4), (253, 172, 3), (251, 173, 1), (253, 183, 1), (253, 195, 4), (251, 195, 1), (254, 191, 1), (255, 193, 3), (254, 194, 1), (255, 194, 1), (255, 193, 1), (255, 194, 1), (251, 184, 1), (253, 172, 1), (255, 171, 1), (254, 170, 0), (252, 176, 34), (254, 168, 94), (254, 150, 70), (255, 142, 56), (252, 139, 44), (253, 137, 44), (253, 135, 45), (252, 132, 38), (252, 129, 22), (250, 124, 7), (248, 121, 0), (249, 119, 1), (251, 118, 1), (249, 117, 0), (248, 115, 0), (248, 114, 0), (248, 115, 0), (248, 114, 1), (248, 114, 1), (248, 114, 0), (249, 113, 0), (249, 113, 0), (248, 112, 1), (247, 110, 1), (249, 112, 3), (249, 111, 4), (250, 111, 2), (250, 111, 1), (250, 112, 1), (250, 112, 0), (250, 112, 1), (249, 113, 1), (249, 113, 0), (249, 113, 0), (250, 114, 0), (250, 114, 1), (252, 115, 3), (252, 115, 3), (252, 115, 3), (252, 115, 1), (252, 115, 1), (253, 117, 2), (253, 117, 2), (253, 117, 2), (252, 116, 2), (252, 116, 1), (253, 117, 0), (253, 117, 1), (253, 117, 2), (253, 117, 2), (253, 117, 1), (253, 118, 0), (255, 119, 1), (254, 120, 1), (254, 121, 1), (253, 122, 1), (253, 124, 1), (253, 123, 1), (254, 124, 2), (254, 126, 2), (254, 127, 1), (253, 129, 1), (254, 131, 1), (254, 132, 2), (253, 133, 1), (254, 136, 1), (251, 137, 17), (252, 141, 39), (253, 144, 53), (254, 145, 64), (253, 146, 67), (255, 157, 83), (111, 61, 44), (117, 73, 11), (213, 131, 3), (203, 129, 2), (207, 135, 6), (220, 67, 11), (225, 4, 2), (227, 0, 1), (225, 1, 1), (226, 0, 1), (226, 0, 1), (226, 0, 1), (227, 1, 2), (227, 1, 2), (227, 1, 2), (227, 1, 2), (227, 1, 2), (226, 0, 1), (226, 0, 1), (214, 80, 2), (214, 77, 2), (212, 72, 0), (213, 72, 1), (216, 71, 0), (219, 72, 2), (222, 70, 3), (220, 63, 3), (218, 50, 1), (212, 44, 0), (235, 94, 21), (248, 130, 33), (232, 111, 2), (231, 102, 0), (232, 97, 0), (232, 93, 0), (232, 92, 0), (233, 92, 0), (232, 92, 0), (231, 91, 0), (229, 89, 0), (224, 85, 1), (220, 82, 1), (215, 78, 0), (216, 81, 0), (193, 61, 9), (126, 2, 4), (123, 0, 0), (119, 0, 0), (166, 70, 40), (255, 218, 112), (254, 196, 72), (253, 187, 40), (255, 182, 13), (255, 181, 3), (254, 179, 1), (252, 179, 0), (253, 180, 0), (253, 180, 0), (252, 180, 0), (253, 182, 0), (255, 184, 1), (253, 187, 0), (253, 190, 1), (253, 190, 0), (252, 194, 0), (253, 198, 2), (253, 200, 8), (252, 201, 11), (252, 202, 8), (254, 198, 5), (253, 178, 2), (250, 155, 1), (254, 152, 1), (255, 155, 1), (255, 155, 1), (252, 154, 0), (252, 171, 7), (254, 191, 7), (254, 195, 2), (254, 197, 3), (254, 198, 2), (254, 196, 2), (254, 193, 5), (251, 177, 4), (250, 158, 0), (254, 164, 2), (255, 170, 4), (254, 171, 0), (253, 175, 43), (254, 161, 87), (254, 145, 63), (255, 139, 53), (253, 134, 35), (251, 134, 28), (252, 132, 37), (252, 129, 31), (250, 126, 13), (248, 123, 1), (248, 119, 0), (249, 117, 0), (250, 116, 1), (248, 114, 0), (247, 113, 1), (248, 113, 1), (248, 113, 1), (248, 113, 1), (248, 112, 1), (249, 112, 1), (248, 111, 1), (248, 111, 1), (248, 111, 2), (247, 110, 1), (248, 111, 3), (248, 111, 2), (249, 111, 0), (249, 110, 0), (250, 110, 0), (250, 110, 0), (250, 111, 0), (249, 112, 2), (249, 112, 0), (249, 112, 1), (248, 112, 1), (249, 112, 1), (249, 112, 2), (249, 112, 2), (250, 113, 2), (251, 114, 3), (251, 114, 3), (252, 115, 2), (252, 115, 2), (251, 115, 1), (252, 115, 2), (252, 115, 2), (252, 116, 1), (252, 116, 1), (252, 116, 2), (253, 116, 1), (253, 117, 1), (253, 117, 1), (254, 118, 2), (254, 118, 0), (253, 118, 0), (252, 120, 0), (252, 122, 0), (254, 123, 1), (255, 125, 2), (254, 126, 2), (254, 126, 1), (253, 127, 2), (252, 129, 1), (253, 131, 1), (253, 132, 2), (254, 132, 0), (251, 132, 6), (253, 137, 32), (255, 140, 45), (254, 140, 51), (252, 141, 51), (255, 157, 79), (122, 73, 45), (108, 67, 8), (211, 130, 4), (206, 128, 2), (206, 133, 3), (210, 116, 7), (214, 21, 4), (228, 0, 5), (224, 0, 1), (226, 0, 1), (226, 0, 1), (226, 0, 1), (227, 1, 2), (227, 1, 2), (227, 1, 2), (227, 1, 2), (227, 1, 2), (226, 0, 1), (226, 0, 1), (205, 76, 1), (205, 71, 1), (208, 71, 1), (211, 71, 0), (215, 68, 1), (215, 64, 2), (214, 61, 0), (224, 71, 3), (231, 79, 8), (221, 80, 16), (238, 111, 29), (232, 106, 8), (224, 94, 1), (224, 91, 0), (225, 88, 0), (226, 85, 0), (226, 85, 0), (224, 85, 2), (224, 85, 2), (225, 84, 2), (224, 83, 2), (220, 80, 0), (215, 77, 0), (211, 73, 1), (209, 69, 0), (204, 72, 3), (144, 23, 5), (118, 0, 1), (115, 0, 0), (190, 108, 53), (255, 210, 79), (255, 182, 32), (253, 177, 7), (253, 176, 0), (253, 173, 1), (252, 170, 2), (252, 170, 2), (254, 171, 2), (254, 172, 1), (254, 173, 0), (254, 175, 1), (254, 177, 2), (255, 179, 1), (255, 181, 1), (255, 182, 1), (255, 184, 2), (255, 186, 2), (254, 188, 0), (254, 189, 1), (255, 188, 0), (254, 186, 0), (251, 178, 3), (252, 153, 1), (255, 143, 0), (255, 143, 0), (254, 143, 0), (253, 144, 0), (252, 150, 1), (252, 163, 1), (252, 175, 5), (253, 180, 6), (254, 179, 6), (253, 174, 4), (251, 164, 2), (250, 155, 1), (251, 153, 2), (252, 157, 0), (254, 163, 3), (254, 169, 0), (253, 170, 51), (252, 151, 77), (255, 139, 54), (254, 134, 47), (252, 131, 29), (250, 130, 21), (250, 127, 29), (248, 124, 17), (249, 124, 2), (248, 121, 1), (247, 118, 1), (249, 115, 0), (248, 113, 0), (248, 113, 1), (247, 112, 2), (247, 111, 2), (247, 111, 3), (246, 111, 3), (248, 111, 3), (248, 110, 3), (247, 110, 2), (247, 110, 2), (247, 110, 2), (247, 110, 1), (248, 110, 1), (248, 110, 0), (247, 110, 1), (247, 110, 2), (249, 109, 0), (249, 109, 0), (249, 110, 1), (248, 110, 3), (248, 110, 3), (248, 110, 3), (248, 110, 3), (248, 110, 2), (248, 111, 2), (248, 110, 1), (249, 111, 2), (250, 112, 4), (250, 112, 4), (250, 113, 2), (250, 113, 1), (250, 113, 2), (251, 114, 3), (251, 114, 3), (251, 114, 2), (251, 114, 1), (251, 114, 1), (252, 115, 0), (252, 115, 0), (252, 115, 0), (252, 116, 2), (253, 116, 0), (252, 117, 0), (252, 119, 0), (253, 120, 0), (255, 121, 0), (255, 123, 0), (254, 125, 0), (254, 124, 0), (254, 125, 1), (253, 127, 0), (254, 128, 0), (254, 129, 2), (254, 130, 1), (253, 130, 1), (252, 132, 12), (253, 133, 26), (254, 136, 43), (253, 137, 44), (255, 151, 70), (132, 78, 46), (84, 48, 10), (204, 125, 10), (204, 126, 2), (203, 126, 3), (202, 128, 3), (208, 88, 9), (216, 8, 5), (226, 0, 2), (226, 0, 2), (224, 0, 1), (226, 0, 0), (227, 0, 0), (226, 0, 0), (227, 0, 0), (229, 0, 0), (228, 0, 0), (226, 0, 0), (226, 0, 0), (195, 68, 1), (199, 67, 1), (203, 67, 1), (205, 66, 0), (205, 59, 0), (212, 63, 3), (235, 85, 8), (250, 105, 5), (255, 123, 7), (255, 129, 24), (231, 105, 14), (218, 90, 1), (219, 84, 3), (217, 80, 0), (219, 80, 0), (220, 80, 1), (220, 79, 2), (220, 79, 4), (220, 79, 2), (219, 79, 1), (218, 78, 2), (214, 77, 1), (210, 74, 1), (207, 70, 1), (205, 67, 2), (203, 70, 2), (159, 39, 6), (116, 0, 1), (114, 0, 0), (209, 128, 57), (255, 197, 41), (255, 173, 2), (252, 171, 0), (251, 169, 1), (252, 167, 1), (252, 165, 3), (252, 164, 2), (252, 164, 1), (254, 165, 1), (254, 166, 1), (254, 169, 0), (254, 170, 0), (253, 171, 1), (254, 174, 1), (254, 176, 1), (253, 178, 1), (255, 180, 2), (255, 181, 3), (255, 181, 4), (255, 180, 3), (254, 178, 2), (253, 174, 1), (253, 151, 2), (254, 139, 1), (254, 141, 1), (254, 141, 0), (254, 145, 1), (255, 151, 3), (254, 153, 0), (253, 153, 0), (253, 153, 0), (254, 155, 0), (253, 154, 0), (252, 153, 0), (253, 154, 0), (252, 152, 1), (252, 151, 0), (251, 153, 1), (251, 157, 0), (252, 162, 52), (251, 145, 71), (254, 134, 47), (252, 131, 33), (249, 129, 15), (249, 127, 18), (248, 124, 21), (248, 121, 11), (248, 120, 1), (248, 118, 2), (247, 116, 1), (248, 114, 0), (248, 111, 1), (247, 111, 0), (247, 110, 1), (246, 109, 2), (245, 109, 3), (246, 109, 3), (247, 110, 3), (247, 110, 3), (246, 108, 2), (246, 108, 2), (246, 108, 2), (247, 108, 2), (249, 109, 3), (249, 109, 2), (249, 109, 2), (249, 109, 3), (249, 109, 3), (249, 109, 2), (249, 109, 3), (249, 109, 2), (249, 108, 3), (249, 109, 3), (249, 109, 3), (249, 109, 3), (249, 109, 2), (248, 108, 1), (248, 108, 2), (249, 109, 3), (249, 109, 3), (249, 110, 2), (249, 110, 1), (250, 111, 2), (250, 111, 2), (250, 111, 2), (250, 112, 1), (249, 113, 1), (250, 112, 1), (251, 112, 0), (251, 112, 0), (250, 113, 1), (252, 114, 1), (254, 115, 0), (253, 117, 1), (253, 117, 1), (255, 119, 0), (255, 120, 1), (255, 121, 1), (253, 122, 0), (253, 122, 0), (255, 123, 1), (255, 124, 0), (255, 125, 0), (253, 126, 1), (254, 127, 2), (254, 128, 1), (252, 128, 1), (252, 129, 11), (254, 134, 31), (253, 134, 36), (255, 141, 41), (144, 82, 42), (50, 32, 13), (179, 111, 11), (207, 124, 1), (201, 120, 1), (197, 118, 0), (199, 122, 4), (198, 86, 5), (210, 11, 0), (218, 0, 0), (216, 0, 3), (218, 14, 15), (222, 31, 28), (222, 37, 33), (224, 38, 34), (225, 30, 26), (220, 13, 7), (216, 8, 5), (224, 14, 10), (186, 56, 4), (190, 56, 1), (191, 53, 0), (187, 45, 0), (190, 44, 3), (226, 82, 7), (242, 99, 4), (243, 100, 0), (241, 103, 0), (237, 103, 0), (215, 89, 1), (209, 80, 1), (210, 77, 0), (210, 75, 0), (211, 74, 1), (213, 75, 2), (213, 75, 3), (213, 76, 1), (213, 75, 1), (212, 74, 0), (210, 72, 1), (205, 72, 0), (202, 70, 0), (201, 67, 1), (199, 64, 1), (199, 67, 3), (167, 45, 12), (112, 0, 0), (114, 2, 3), (220, 134, 56), (255, 187, 18), (253, 171, 0), (251, 168, 0), (251, 163, 0), (250, 162, 0), (250, 161, 0), (251, 161, 1), (251, 161, 0), (251, 161, 0), (253, 161, 0), (254, 162, 0), (253, 164, 1), (253, 166, 1), (253, 169, 0), (254, 171, 0), (253, 173, 0), (254, 175, 1), (254, 176, 1), (254, 177, 1), (254, 177, 1), (254, 175, 0), (252, 169, 0), (252, 148, 2), (254, 134, 3), (254, 137, 1), (252, 138, 1), (253, 142, 1), (255, 149, 3), (255, 151, 1), (254, 151, 0), (253, 152, 0), (254, 153, 0), (255, 153, 0), (255, 153, 0), (255, 153, 0), (254, 151, 0), (252, 147, 0), (252, 148, 0), (251, 152, 0), (252, 158, 55), (252, 144, 68), (252, 132, 34), (250, 129, 14), (247, 125, 3), (247, 123, 7), (248, 122, 7), (247, 118, 2), (248, 118, 2), (248, 117, 2), (246, 115, 0), (245, 114, 0), (246, 111, 1), (245, 110, 1), (244, 109, 2), (245, 108, 3), (246, 108, 1), (247, 108, 2), (246, 108, 2), (246, 108, 2), (246, 108, 2), (246, 108, 2), (248, 108, 2), (248, 107, 2), (247, 108, 2), (248, 109, 2), (249, 109, 1), (248, 108, 1), (248, 107, 3), (248, 108, 2), (248, 108, 1), (247, 107, 2), (247, 107, 2), (248, 108, 2), (248, 108, 2), (248, 108, 2), (248, 108, 2), (247, 107, 1), (246, 106, 1), (246, 106, 1), (245, 106, 1), (246, 108, 0), (247, 108, 0), (247, 109, 1), (248, 110, 2), (249, 110, 2), (249, 111, 2), (248, 111, 2), (249, 111, 2), (251, 111, 2), (252, 110, 2), (251, 111, 2), (252, 113, 1), (253, 114, 1), (253, 115, 0), (252, 116, 0), (253, 117, 0), (254, 118, 1), (255, 118, 1), (254, 118, 1), (253, 119, 0), (253, 120, 1), (255, 121, 1), (255, 122, 0), (253, 123, 1), (253, 124, 0), (253, 125, 0), (253, 124, 0), (253, 125, 2), (253, 127, 7), (253, 125, 10), (255, 134, 28), (149, 83, 37), (34, 25, 10), (124, 75, 14), (205, 123, 5), (193, 116, 0), (188, 111, 0), (184, 106, 0), (188, 116, 11), (209, 115, 54), (228, 110, 93), (241, 131, 129), (245, 147, 138), (251, 158, 148), (251, 160, 151), (251, 161, 153), (250, 156, 146), (244, 138, 126), (245, 134, 125), (252, 138, 129), (183, 48, 7), (186, 48, 2), (184, 43, 2), (178, 34, 1), (194, 49, 8), (228, 88, 6), (233, 92, 0), (233, 90, 0), (230, 86, 1), (222, 82, 1), (207, 78, 3), (205, 73, 1), (205, 72, 0), (204, 70, 0), (205, 70, 0), (206, 70, 1), (206, 70, 2), (207, 70, 2), (206, 70, 1), (205, 70, 1), (203, 68, 1), (200, 67, 1), (199, 65, 1), (197, 62, 1), (192, 60, 1), (193, 63, 5), (166, 43, 12), (109, 0, 3), (118, 10, 21), (199, 109, 37), (255, 183, 13), (251, 168, 0), (250, 165, 0), (250, 160, 0), (250, 158, 0), (250, 157, 0), (250, 158, 0), (250, 158, 0), (251, 158, 0), (253, 157, 0), (253, 158, 0), (253, 160, 1), (253, 162, 1), (253, 164, 0), (254, 167, 0), (254, 169, 0), (255, 171, 2), (254, 173, 2), (254, 174, 1), (255, 174, 1), (254, 172, 0), (251, 166, 0), (252, 142, 0), (253, 125, 0), (252, 126, 0), (249, 128, 0), (250, 134, 0), (253, 142, 0), (252, 144, 0), (252, 144, 0), (253, 146, 0), (252, 149, 0), (254, 152, 1), (255, 154, 1), (255, 153, 2), (255, 149, 0), (253, 145, 0), (254, 148, 1), (251, 156, 3), (250, 157, 55), (250, 139, 62), (250, 129, 26), (250, 126, 5), (249, 123, 1), (249, 120, 1), (247, 117, 0), (246, 115, 1), (247, 114, 2), (248, 114, 2), (247, 114, 1), (247, 113, 2), (246, 110, 3), (245, 109, 2), (245, 109, 1), (246, 108, 3), (246, 107, 1), (247, 107, 1), (246, 107, 1), (245, 107, 1), (246, 107, 1), (246, 107, 1), (247, 107, 1), (247, 106, 1), (246, 107, 1), (246, 107, 1), (246, 106, 0), (247, 107, 1), (247, 106, 2), (247, 107, 1), (247, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (247, 107, 1), (247, 107, 1), (248, 107, 2), (248, 106, 1), (248, 106, 1), (248, 107, 2), (248, 107, 2), (247, 107, 1), (248, 107, 1), (248, 107, 1), (249, 107, 2), (249, 108, 2), (248, 109, 2), (248, 109, 2), (248, 109, 2), (248, 110, 2), (249, 110, 2), (249, 110, 1), (250, 111, 1), (252, 113, 2), (252, 113, 2), (251, 114, 1), (253, 114, 1), (254, 114, 2), (255, 114, 2), (254, 115, 0), (252, 116, 0), (252, 118, 1), (253, 120, 2), (254, 120, 1), (254, 120, 1), (254, 122, 1), (254, 122, 1), (254, 122, 1), (253, 121, 1), (252, 121, 1), (252, 119, 1), (255, 131, 30), (145, 80, 38), (37, 27, 16), (58, 35, 15), (158, 101, 12), (184, 107, 0), (187, 107, 18), (217, 137, 73), (244, 162, 138), (252, 170, 169), (254, 161, 161), (255, 144, 133), (254, 137, 121), (251, 132, 116), (251, 130, 118), (252, 130, 123), (253, 133, 128), (253, 140, 132), (255, 142, 136), (254, 145, 143), (181, 42, 4), (186, 47, 3), (183, 41, 1), (177, 34, 0), (188, 47, 5), (225, 84, 6), (227, 85, 1), (226, 83, 3), (223, 79, 0), (217, 74, 0), (203, 72, 1), (202, 70, 1), (201, 68, 0), (200, 67, 0), (200, 67, 0), (200, 67, 1), (200, 67, 1), (199, 66, 1), (199, 66, 0), (199, 66, 0), (199, 65, 1), (197, 63, 1), (196, 60, 1), (192, 58, 2), (187, 57, 1), (186, 58, 5), (152, 33, 7), (113, 7, 9), (117, 5, 18), (165, 65, 5), (255, 179, 10), (252, 167, 0), (250, 163, 1), (249, 159, 0), (250, 157, 0), (250, 155, 0), (249, 154, 0), (248, 154, 0), (250, 155, 0), (252, 155, 1), (252, 155, 1), (252, 156, 0), (253, 159, 0), (253, 160, 0), (254, 162, 0), (255, 165, 1), (255, 168, 1), (255, 170, 1), (254, 172, 1), (255, 171, 1), (254, 168, 0), (251, 154, 0), (248, 133, 0), (246, 142, 16), (246, 171, 42), (249, 187, 58), (250, 195, 60), (251, 196, 51), (250, 188, 34), (248, 178, 19), (249, 164, 6), (251, 152, 0), (251, 148, 0), (254, 150, 0), (255, 152, 3), (255, 147, 1), (254, 147, 1), (253, 156, 3), (253, 167, 7), (250, 160, 56), (248, 133, 54), (250, 126, 21), (249, 125, 10), (249, 120, 1), (248, 117, 2), (247, 114, 2), (246, 112, 1), (248, 112, 1), (247, 112, 1), (248, 112, 2), (248, 111, 3), (247, 110, 3), (246, 109, 2), (246, 108, 2), (246, 108, 2), (245, 107, 1), (245, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (245, 106, 1), (245, 106, 0), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (248, 108, 2), (248, 106, 1), (248, 106, 1), (249, 107, 2), (249, 107, 2), (249, 107, 2), (249, 107, 2), (249, 106, 2), (249, 106, 2), (248, 107, 2), (247, 107, 2), (247, 107, 2), (247, 107, 2), (247, 110, 1), (247, 110, 1), (247, 110, 1), (250, 111, 1), (251, 112, 2), (252, 112, 3), (253, 112, 2), (252, 112, 3), (253, 113, 1), (253, 113, 1), (251, 113, 1), (251, 115, 0), (252, 115, 0), (253, 117, 2), (254, 118, 1), (254, 118, 0), (255, 119, 1), (255, 119, 1), (254, 119, 1), (252, 118, 0), (253, 118, 0), (252, 117, 0), (255, 127, 31), (139, 75, 39), (44, 28, 18), (38, 27, 17), (80, 39, 13), (202, 123, 68), (246, 154, 137), (255, 154, 160), (255, 141, 140), (253, 118, 109), (249, 105, 91), (252, 101, 81), (254, 100, 84), (252, 98, 86), (252, 97, 88), (253, 98, 91), (254, 101, 94), (252, 104, 98), (252, 107, 102), (252, 113, 109), (174, 42, 1), (172, 39, 2), (169, 33, 1), (163, 25, 1), (157, 18, 2), (195, 59, 9), (227, 86, 6), (226, 84, 1), (222, 79, 0), (221, 77, 0), (208, 73, 1), (199, 67, 2), (197, 66, 2), (196, 66, 0), (196, 66, 0), (196, 65, 1), (196, 66, 0), (195, 64, 0), (195, 64, 0), (197, 64, 1), (197, 64, 1), (195, 61, 1), (194, 59, 2), (190, 57, 2), (184, 55, 2), (182, 52, 4), (131, 11, 0), (121, 12, 11), (114, 9, 14), (139, 59, 41), (248, 167, 23), (255, 166, 0), (251, 163, 4), (249, 158, 0), (250, 157, 0), (250, 154, 0), (250, 153, 1), (248, 153, 1), (248, 152, 1), (250, 151, 2), (249, 151, 1), (249, 152, 0), (251, 154, 0), (253, 156, 1), (253, 159, 0), (254, 163, 1), (255, 166, 0), (254, 169, 1), (254, 172, 3), (254, 166, 0), (249, 158, 0), (248, 172, 41), (249, 208, 101), (250, 236, 142), (253, 245, 152), (255, 243, 147), (255, 241, 138), (254, 237, 124), (255, 232, 106), (252, 228, 92), (253, 219, 80), (252, 208, 55), (247, 188, 30), (251, 158, 6), (252, 141, 0), (253, 144, 0), (252, 153, 3), (251, 164, 2), (254, 174, 5), (253, 161, 57), (249, 129, 55), (249, 124, 24), (248, 127, 32), (249, 120, 7), (246, 116, 2), (246, 113, 2), (247, 110, 0), (247, 110, 1), (246, 111, 1), (247, 110, 2), (247, 109, 2), (247, 110, 2), (246, 109, 3), (246, 108, 3), (246, 108, 2), (245, 107, 1), (245, 107, 1), (246, 106, 1), (247, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 107, 1), (244, 107, 0), (244, 106, 0), (245, 107, 2), (246, 106, 2), (247, 106, 1), (248, 106, 1), (248, 108, 2), (247, 107, 1), (247, 105, 1), (247, 105, 1), (247, 106, 1), (248, 106, 1), (248, 106, 1), (248, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (247, 106, 1), (246, 106, 1), (247, 108, 1), (248, 109, 1), (249, 109, 1), (250, 111, 1), (251, 111, 1), (252, 110, 3), (252, 111, 4), (251, 112, 2), (251, 112, 1), (251, 112, 1), (251, 112, 2), (250, 112, 0), (251, 112, 0), (253, 113, 1), (253, 114, 2), (252, 116, 0), (254, 116, 1), (255, 116, 1), (254, 116, 1), (253, 116, 0), (253, 115, 0), (254, 114, 0), (255, 123, 29), (129, 66, 35), (34, 24, 10), (77, 39, 23), (189, 106, 101), (255, 143, 143), (255, 124, 124), (254, 109, 110), (255, 94, 82), (254, 81, 67), (253, 79, 65), (254, 78, 62), (255, 77, 63), (255, 75, 65), (255, 76, 66), (255, 75, 66), (254, 76, 69), (251, 79, 73), (251, 84, 77), (252, 88, 82), (172, 52, 3), (167, 46, 4), (165, 41, 1), (160, 30, 6), (135, 13, 3), (142, 30, 2), (196, 66, 9), (215, 77, 5), (215, 79, 7), (205, 67, 10), (191, 55, 3), (197, 64, 0), (197, 65, 1), (196, 65, 1), (195, 64, 0), (194, 63, 1), (194, 63, 0), (194, 64, 1), (197, 63, 1), (197, 64, 2), (195, 62, 1), (192, 60, 0), (189, 58, 1), (187, 56, 3), (185, 47, 0), (158, 34, 0), (133, 68, 68), (161, 150, 165), (170, 188, 203), (179, 217, 237), (222, 188, 110), (253, 162, 0), (251, 163, 3), (251, 158, 1), (250, 155, 2), (249, 154, 2), (249, 153, 2), (247, 151, 0), (247, 149, 0), (247, 148, 1), (245, 148, 0), (246, 150, 0), (249, 153, 0), (253, 155, 1), (254, 158, 0), (254, 162, 1), (255, 164, 3), (255, 165, 2), (253, 159, 0), (243, 164, 12), (248, 206, 92), (252, 240, 149), (251, 246, 154), (252, 239, 146), (254, 236, 140), (252, 234, 134), (252, 235, 126), (254, 234, 124), (255, 232, 121), (255, 231, 118), (255, 230, 113), (253, 231, 107), (252, 232, 105), (252, 218, 92), (247, 178, 41), (247, 145, 0), (252, 154, 0), (252, 166, 1), (253, 178, 4), (253, 170, 60), (248, 133, 62), (249, 123, 23), (246, 122, 22), (246, 117, 7), (245, 115, 4), (246, 111, 1), (246, 108, 0), (245, 109, 2), (244, 109, 2), (244, 109, 2), (245, 108, 2), (246, 108, 2), (246, 108, 2), (246, 108, 2), (246, 108, 2), (245, 107, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (245, 105, 0), (243, 106, 0), (243, 106, 0), (244, 106, 1), (245, 107, 3), (246, 106, 2), (248, 106, 1), (249, 105, 1), (248, 106, 1), (247, 105, 0), (246, 104, 0), (246, 104, 0), (245, 105, 0), (247, 106, 1), (248, 106, 1), (248, 106, 1), (246, 106, 1), (246, 106, 1), (248, 106, 1), (248, 106, 1), (246, 106, 1), (247, 107, 2), (249, 108, 3), (251, 108, 3), (251, 109, 3), (251, 109, 3), (250, 110, 4), (249, 109, 3), (250, 109, 1), (251, 110, 1), (251, 110, 2), (251, 110, 3), (251, 110, 1), (251, 110, 1), (252, 110, 2), (252, 111, 2), (251, 113, 1), (253, 113, 2), (254, 113, 2), (254, 113, 2), (254, 113, 2), (254, 112, 1), (255, 110, 0), (249, 118, 26), (88, 47, 16), (78, 41, 33), (219, 116, 104), (255, 121, 115), (249, 103, 103), (247, 92, 89), (250, 80, 77), (251, 65, 51), (254, 61, 46), (252, 60, 45), (250, 58, 42), (251, 58, 43), (251, 57, 44), (250, 58, 46), (252, 60, 50), (251, 61, 53), (249, 64, 57), (250, 67, 61), (251, 70, 66), (164, 51, 2), (160, 49, 3), (158, 45, 2), (154, 38, 2), (157, 43, 5), (164, 52, 4), (164, 45, 1), (168, 46, 1), (169, 46, 5), (147, 22, 5), (134, 21, 1), (159, 49, 4), (192, 70, 6), (199, 66, 1), (195, 64, 2), (194, 64, 1), (194, 63, 1), (195, 65, 2), (195, 64, 2), (195, 63, 2), (193, 61, 1), (187, 59, 1), (186, 57, 2), (180, 46, 0), (165, 68, 26), (165, 160, 149), (165, 223, 240), (169, 234, 255), (169, 232, 253), (174, 229, 255), (185, 211, 214), (240, 168, 36), (253, 158, 0), (242, 154, 1), (243, 153, 1), (247, 154, 1), (248, 153, 1), (248, 153, 1), (248, 151, 0), (247, 149, 0), (244, 149, 0), (245, 151, 0), (249, 153, 1), (252, 154, 2), (253, 155, 0), (253, 158, 1), (255, 160, 1), (252, 153, 0), (243, 161, 13), (252, 213, 102), (254, 239, 152), (250, 235, 127), (251, 232, 113), (252, 230, 110), (253, 230, 106), (252, 230, 104), (252, 228, 104), (253, 228, 106), (254, 230, 104), (253, 229, 104), (252, 230, 109), (253, 231, 121), (252, 232, 131), (254, 234, 140), (255, 236, 137), (248, 202, 67), (246, 159, 1), (252, 160, 0), (253, 190, 3), (248, 180, 51), (245, 136, 77), (246, 124, 31), (244, 119, 5), (243, 116, 2), (245, 113, 3), (246, 111, 1), (246, 109, 0), (246, 109, 1), (245, 108, 1), (245, 107, 1), (245, 107, 1), (246, 108, 2), (246, 108, 2), (246, 108, 2), (246, 108, 2), (245, 107, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (244, 106, 0), (244, 106, 0), (244, 106, 0), (244, 106, 0), (244, 106, 0), (244, 105, 1), (242, 104, 2), (244, 106, 1), (245, 105, 0), (246, 105, 0), (246, 105, 0), (247, 105, 0), (244, 105, 0), (243, 105, 0), (244, 104, 0), (244, 104, 0), (244, 105, 0), (244, 104, 0), (245, 104, 0), (244, 104, 0), (244, 104, 0), (244, 104, 0), (245, 105, 0), (246, 106, 1), (247, 107, 2), (248, 108, 3), (249, 108, 3), (250, 108, 2), (250, 108, 3), (250, 108, 3), (250, 108, 3), (249, 108, 1), (250, 108, 1), (250, 108, 2), (250, 108, 3), (249, 107, 2), (249, 107, 1), (250, 108, 2), (251, 108, 1), (252, 109, 1), (253, 110, 2), (252, 111, 2), (254, 110, 2), (255, 109, 3), (254, 109, 2), (255, 106, 0), (227, 98, 26), (126, 54, 37), (221, 106, 100), (255, 101, 98), (247, 85, 80), (243, 82, 77), (241, 74, 72), (247, 63, 53), (246, 53, 29), (248, 50, 25), (248, 48, 24), (246, 45, 22), (245, 47, 25), (247, 49, 31), (243, 47, 29), (244, 48, 33), (245, 50, 38), (244, 53, 45), (244, 54, 49), (241, 58, 53), (156, 51, 3), (153, 48, 3), (148, 42, 0), (150, 43, 2), (164, 60, 2), (162, 54, 1), (152, 44, 0), (145, 38, 0), (142, 29, 0), (135, 27, 4), (116, 43, 33), (104, 41, 45), (131, 44, 18), (184, 64, 7), (197, 68, 7), (196, 65, 3), (193, 64, 1), (193, 64, 2), (193, 64, 4), (192, 63, 2), (190, 60, 1), (183, 59, 2), (183, 46, 0), (174, 70, 35), (167, 190, 190), (141, 221, 255), (131, 199, 242), (128, 185, 233), (110, 172, 237), (100, 157, 235), (92, 150, 245), (152, 146, 169), (244, 158, 12), (245, 153, 0), (241, 152, 3), (247, 155, 1), (251, 156, 2), (251, 156, 2), (251, 153, 1), (249, 150, 1), (247, 150, 2), (246, 150, 1), (248, 150, 0), (250, 151, 0), (253, 153, 1), (254, 154, 2), (253, 150, 0), (247, 151, 7), (250, 207, 77), (255, 230, 121), (254, 225, 97), (254, 224, 85), (255, 222, 83), (255, 222, 77), (255, 223, 76), (254, 223, 77), (254, 222, 77), (254, 222, 79), (253, 223, 82), (252, 225, 88), (252, 227, 101), (254, 230, 116), (254, 231, 127), (255, 232, 137), (255, 233, 150), (255, 238, 148), (248, 206, 66), (250, 161, 0), (255, 193, 3), (251, 179, 32), (245, 138, 80), (244, 125, 41), (245, 118, 7), (243, 117, 1), (244, 114, 2), (245, 110, 2), (245, 108, 2), (246, 107, 1), (245, 106, 0), (244, 106, 0), (244, 106, 0), (245, 107, 1), (245, 107, 1), (245, 107, 1), (245, 107, 1), (245, 107, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (246, 106, 1), (245, 106, 0), (244, 106, 2), (244, 106, 2), (242, 105, 1), (243, 105, 1), (243, 104, 1), (242, 104, 1), (242, 105, 1), (243, 104, 1), (243, 104, 1), (243, 104, 1), (244, 104, 1), (243, 104, 1), (244, 104, 1), (246, 103, 1), (245, 104, 1), (244, 103, 0), (244, 102, 0), (244, 102, 0), (244, 102, 0), (245, 103, 1), (245, 103, 1), (246, 104, 1), (246, 104, 1), (247, 105, 2), (247, 105, 2), (247, 106, 1), (249, 107, 1), (249, 107, 2), (249, 107, 2), (249, 107, 1), (249, 107, 1), (249, 107, 1), (249, 107, 1), (249, 107, 2), (249, 107, 2), (249, 107, 2), (249, 106, 2), (251, 106, 2), (251, 106, 0), (252, 108, 1), (251, 107, 1), (252, 106, 2), (254, 105, 2), (255, 105, 2), (253, 101, 0), (245, 98, 34), (243, 90, 85), (249, 80, 71), (238, 68, 61), (238, 68, 61), (235, 65, 57), (238, 60, 52), (242, 45, 27), (242, 39, 15), (242, 37, 11), (243, 34, 10), (242, 32, 8), (240, 38, 14), (243, 38, 17), (239, 31, 12), (242, 36, 14), (241, 37, 19), (239, 39, 27), (239, 42, 36), (237, 48, 41), (137, 47, 0), (133, 45, 0), (129, 37, 0), (143, 43, 1), (157, 55, 0), (150, 59, 11), (156, 74, 49), (161, 80, 64), (147, 55, 40), (117, 35, 24), (102, 55, 68), (88, 53, 70), (79, 25, 43), (100, 31, 21), (151, 50, 8), (182, 63, 6), (191, 66, 8), (195, 67, 7), (194, 67, 3), (191, 65, 2), (187, 64, 2), (174, 52, 0), (141, 51, 10), (149, 173, 178), (120, 198, 245), (88, 169, 232), (63, 152, 236), (38, 131, 229), (15, 119, 229), (4, 119, 236), (5, 119, 238), (18, 119, 245), (128, 135, 155), (244, 153, 20), (250, 150, 0), (246, 153, 3), (249, 155, 1), (248, 153, 1), (248, 152, 0), (247, 150, 1), (246, 148, 2), (245, 148, 1), (247, 149, 0), (247, 148, 0), (250, 149, 2), (250, 147, 0), (246, 141, 0), (250, 184, 49), (254, 221, 95), (252, 217, 86), (251, 217, 63), (251, 215, 56), (252, 214, 55), (253, 214, 52), (254, 214, 53), (255, 213, 54), (254, 213, 55), (254, 215, 56), (253, 216, 63), (253, 218, 76), (254, 220, 89), (254, 223, 105), (253, 227, 116), (254, 230, 129), (255, 232, 141), (255, 235, 151), (253, 235, 120), (248, 183, 20), (251, 185, 0), (249, 186, 37), (241, 141, 75), (246, 128, 53), (245, 119, 14), (243, 114, 1), (244, 113, 3), (244, 111, 2), (245, 109, 2), (245, 108, 1), (244, 106, 0), (244, 106, 0), (244, 106, 0), (245, 107, 1), (245, 107, 1), (245, 107, 1), (245, 107, 1), (245, 107, 1), (245, 106, 0), (245, 106, 0), (245, 106, 0), (245, 106, 0), (245, 106, 0), (245, 106, 0), (245, 106, 0), (244, 107, 1), (243, 105, 1), (243, 105, 2), (243, 105, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (244, 104, 1), (245, 102, 0), (245, 102, 0), (244, 102, 0), (244, 102, 0), (244, 102, 0), (244, 102, 0), (246, 103, 1), (246, 103, 1), (246, 103, 1), (246, 103, 1), (246, 103, 2), (246, 103, 2), (246, 104, 1), (248, 105, 1), (248, 105, 1), (248, 105, 1), (247, 105, 1), (248, 106, 1), (248, 106, 1), (248, 106, 1), (248, 106, 1), (247, 104, 0), (247, 104, 0), (248, 104, 0), (248, 104, 0), (249, 104, 0), (251, 105, 0), (251, 104, 0), (252, 102, 1), (254, 101, 2), (253, 97, 1), (249, 94, 3), (250, 83, 34), (243, 56, 36), (239, 45, 19), (237, 44, 24), (235, 48, 28), (234, 53, 38), (231, 46, 26), (233, 29, 2), (234, 26, 2), (233, 23, 0), (237, 22, 0), (238, 21, 0), (235, 24, 3), (238, 21, 3), (235, 15, 1), (236, 17, 1), (236, 20, 3), (236, 24, 9), (239, 28, 16), (238, 34, 29), (123, 36, 0), (120, 35, 0), (116, 30, 1), (127, 30, 0), (129, 52, 28), (144, 117, 140), (152, 147, 201), (165, 149, 208), (187, 141, 184), (152, 97, 125), (88, 50, 62), (79, 43, 54), (77, 35, 47), (76, 30, 35), (78, 26, 21), (86, 23, 8), (105, 27, 10), (117, 38, 12), (123, 40, 7), (121, 35, 11), (105, 30, 9), (80, 16, 1), (112, 107, 110), (99, 184, 247), (46, 151, 237), (31, 147, 234), (6, 127, 234), (0, 113, 230), (0, 111, 230), (0, 110, 233), (1, 109, 231), (0, 109, 228), (0, 110, 235), (92, 120, 167), (208, 142, 44), (246, 149, 0), (247, 152, 0), (244, 149, 0), (244, 148, 1), (242, 146, 3), (241, 146, 3), (242, 145, 2), (243, 145, 1), (242, 144, 1), (244, 142, 0), (242, 134, 0), (241, 153, 13), (255, 202, 63), (255, 206, 69), (254, 206, 54), (253, 205, 31), (255, 203, 23), (255, 201, 21), (254, 202, 19), (254, 203, 19), (254, 202, 19), (254, 202, 20), (254, 204, 28), (255, 207, 47), (255, 210, 65), (255, 212, 77), (254, 215, 91), (252, 222, 98), (252, 227, 113), (253, 230, 128), (253, 234, 138), (254, 235, 129), (247, 208, 59), (249, 221, 75), (250, 234, 122), (239, 145, 71), (244, 126, 56), (242, 121, 24), (245, 114, 4), (246, 112, 1), (243, 110, 1), (244, 109, 1), (244, 108, 1), (244, 106, 1), (244, 106, 0), (244, 105, 1), (245, 107, 1), (245, 107, 1), (245, 107, 1), (245, 107, 1), (245, 107, 1), (246, 106, 0), (244, 106, 0), (243, 106, 0), (243, 106, 0), (243, 106, 0), (244, 106, 1), (244, 106, 0), (242, 106, 1), (242, 105, 2), (242, 104, 1), (242, 105, 0), (242, 104, 1), (242, 104, 1), (242, 104, 1), (244, 104, 1), (244, 104, 1), (243, 104, 1), (243, 104, 1), (242, 104, 2), (242, 103, 1), (242, 103, 1), (242, 103, 1), (244, 102, 0), (245, 101, 0), (245, 102, 0), (244, 102, 0), (244, 102, 0), (244, 102, 0), (246, 103, 1), (246, 103, 1), (246, 103, 1), (246, 103, 1), (246, 102, 1), (246, 103, 1), (246, 102, 1), (246, 102, 1), (246, 102, 1), (246, 103, 1), (246, 103, 1), (247, 103, 1), (247, 104, 1), (248, 105, 1), (248, 105, 1), (247, 104, 0), (247, 104, 0), (247, 103, 0), (247, 101, 0), (248, 101, 0), (249, 102, 1), (250, 101, 0), (251, 99, 2), (252, 96, 3), (252, 88, 1), (245, 71, 2), (232, 42, 12), (231, 28, 2), (230, 22, 0), (231, 20, 3), (230, 19, 4), (230, 24, 17), (227, 17, 15), (228, 3, 0), (230, 4, 2), (228, 3, 1), (230, 4, 2), (231, 5, 2), (228, 5, 1), (231, 10, 4), (228, 8, 2), (225, 5, 0), (227, 9, 2), (228, 11, 4), (228, 16, 5), (230, 24, 19), (112, 27, 8), (112, 25, 10), (109, 18, 0), (114, 23, 1), (131, 96, 135), (108, 123, 190), (95, 121, 184), (97, 122, 187), (136, 122, 181), (154, 108, 149), (108, 64, 79), (69, 28, 39), (75, 34, 42), (80, 35, 40), (76, 30, 37), (50, 6, 27), (37, 2, 27), (34, 2, 21), (32, 4, 19), (29, 5, 20), (31, 0, 10), (46, 19, 41), (69, 140, 206), (16, 140, 234), (0, 135, 229), (3, 129, 229), (2, 107, 221), (1, 101, 223), (1, 100, 226), (1, 96, 225), (2, 96, 223), (1, 97, 220), (0, 100, 218), (0, 98, 231), (36, 104, 187), (127, 119, 103), (207, 133, 35), (235, 140, 0), (240, 140, 0), (239, 139, 0), (235, 143, 2), (236, 141, 2), (237, 140, 1), (243, 141, 5), (238, 136, 5), (229, 126, 1), (243, 171, 33), (248, 198, 52), (252, 196, 38), (253, 194, 23), (251, 194, 8), (252, 193, 3), (253, 192, 2), (252, 192, 1), (252, 192, 1), (253, 192, 1), (252, 193, 0), (253, 196, 8), (254, 199, 38), (254, 201, 59), (254, 204, 65), (253, 210, 68), (254, 214, 79), (254, 218, 94), (253, 224, 101), (254, 229, 110), (254, 231, 113), (254, 234, 101), (253, 238, 99), (254, 235, 80), (241, 155, 63), (237, 120, 54), (242, 123, 36), (246, 114, 14), (245, 110, 1), (242, 109, 1), (244, 107, 1), (244, 106, 0), (243, 105, 0), (242, 104, 1), (242, 104, 1), (244, 106, 0), (244, 106, 0), (244, 107, 0), (246, 107, 1), (246, 106, 1), (247, 106, 1), (245, 107, 1), (243, 107, 0), (242, 105, 0), (243, 105, 2), (244, 106, 2), (244, 106, 2), (244, 106, 2), (243, 105, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (241, 103, 0), (243, 103, 0), (245, 103, 1), (245, 103, 1), (244, 104, 1), (243, 103, 2), (243, 102, 2), (242, 101, 0), (242, 101, 0), (243, 101, 1), (244, 101, 2), (244, 101, 2), (244, 102, 0), (244, 102, 0), (244, 102, 0), (244, 102, 0), (244, 102, 0), (245, 102, 0), (247, 102, 2), (247, 102, 1), (247, 101, 0), (246, 101, 0), (246, 100, 1), (246, 100, 2), (246, 100, 1), (246, 101, 0), (246, 101, 1), (246, 101, 1), (247, 102, 1), (247, 102, 1), (246, 102, 1), (245, 102, 1), (247, 101, 2), (247, 100, 2), (247, 99, 2), (247, 99, 2), (246, 100, 0), (248, 99, 1), (249, 95, 3), (248, 90, 3), (249, 76, 6), (230, 34, 0), (222, 10, 1), (222, 8, 1), (222, 4, 0), (224, 4, 0), (222, 2, 0), (221, 0, 0), (225, 1, 2), (225, 0, 2), (226, 0, 3), (227, 0, 1), (224, 0, 0), (224, 0, 0), (223, 0, 1), (224, 2, 4), (223, 3, 2), (222, 2, 0), (221, 1, 0), (221, 0, 1), (218, 3, 4), (222, 13, 14), (113, 50, 133), (114, 47, 139), (105, 35, 100), (102, 38, 70), (95, 63, 121), (74, 53, 121), (76, 54, 131), (68, 78, 144), (78, 89, 142), (103, 78, 112), (105, 58, 74), (70, 23, 35), (67, 26, 37), (72, 32, 41), (61, 23, 34), (43, 9, 36), (39, 11, 39), (40, 14, 36), (35, 15, 36), (30, 12, 30), (29, 12, 25), (41, 91, 154), (7, 126, 233), (0, 118, 220), (3, 112, 218), (2, 105, 214), (0, 95, 206), (1, 91, 207), (1, 90, 209), (0, 88, 210), (1, 87, 211), (1, 88, 207), (1, 88, 204), (1, 91, 206), (0, 91, 211), (0, 90, 210), (29, 95, 182), (89, 106, 125), (140, 115, 85), (179, 121, 57), (184, 111, 13), (192, 113, 13), (181, 109, 12), (153, 88, 12), (156, 96, 28), (224, 159, 50), (241, 179, 35), (246, 188, 28), (246, 189, 11), (246, 187, 1), (246, 185, 1), (246, 184, 1), (247, 183, 1), (248, 183, 0), (250, 183, 0), (251, 182, 0), (252, 183, 1), (253, 186, 1), (253, 188, 15), (253, 191, 36), (252, 196, 45), (251, 201, 51), (254, 205, 60), (255, 209, 66), (254, 216, 60), (255, 221, 63), (254, 224, 62), (250, 219, 34), (248, 212, 11), (255, 213, 6), (246, 171, 30), (235, 119, 60), (242, 119, 43), (243, 115, 12), (243, 109, 1), (242, 108, 1), (242, 107, 0), (241, 106, 0), (242, 104, 1), (242, 104, 1), (242, 105, 0), (244, 106, 0), (244, 106, 0), (244, 106, 0), (244, 106, 0), (244, 106, 0), (244, 107, 1), (244, 107, 1), (244, 106, 1), (242, 104, 2), (243, 105, 1), (244, 106, 1), (244, 106, 2), (244, 106, 2), (243, 105, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 103, 0), (243, 103, 0), (244, 102, 0), (244, 102, 0), (243, 103, 0), (242, 102, 0), (242, 101, 0), (242, 101, 0), (242, 101, 0), (243, 101, 1), (244, 101, 2), (244, 101, 2), (244, 102, 0), (244, 102, 0), (244, 102, 0), (244, 102, 0), (244, 102, 0), (246, 100, 2), (246, 100, 3), (246, 101, 3), (244, 100, 1), (245, 99, 0), (245, 99, 0), (246, 100, 2), (246, 100, 2), (246, 100, 2), (246, 100, 2), (246, 100, 2), (245, 100, 0), (245, 100, 0), (245, 100, 1), (245, 100, 2), (247, 99, 2), (247, 98, 2), (246, 98, 2), (246, 98, 2), (246, 97, 1), (247, 94, 2), (246, 89, 0), (245, 83, 4), (239, 53, 8), (218, 5, 0), (217, 0, 2), (217, 1, 3), (220, 1, 1), (221, 2, 0), (220, 1, 0), (219, 0, 0), (221, 1, 0), (220, 0, 0), (220, 0, 1), (220, 0, 0), (219, 1, 0), (217, 1, 0), (219, 1, 0), (219, 0, 1), (218, 1, 1), (216, 1, 0), (216, 0, 0), (216, 0, 2), (215, 1, 4), (214, 4, 12), (76, 28, 147), (74, 29, 145), (71, 30, 143), (80, 34, 136), (64, 14, 91), (53, 0, 66), (61, 0, 74), (71, 6, 82), (69, 50, 105), (74, 72, 102), (91, 56, 69), (72, 18, 20), (44, 3, 8), (33, 6, 14), (22, 3, 8), (33, 13, 36), (42, 16, 46), (42, 18, 42), (34, 15, 37), (34, 7, 24), (38, 63, 106), (10, 126, 220), (1, 107, 215), (1, 102, 206), (2, 93, 206), (2, 88, 202), (0, 88, 200), (0, 85, 198), (0, 81, 196), (0, 79, 195), (1, 80, 194), (0, 79, 190), (0, 78, 186), (1, 77, 192), (1, 79, 189), (0, 80, 186), (0, 82, 195), (0, 86, 205), (0, 93, 209), (34, 104, 202), (51, 55, 95), (37, 18, 11), (28, 21, 12), (11, 4, 11), (95, 58, 40), (225, 164, 49), (239, 176, 16), (242, 180, 3), (241, 181, 0), (241, 179, 0), (241, 178, 0), (243, 177, 1), (245, 176, 2), (246, 176, 1), (247, 175, 0), (248, 174, 0), (249, 175, 0), (250, 176, 0), (250, 178, 2), (252, 181, 7), (252, 184, 12), (251, 190, 18), (254, 193, 26), (253, 196, 29), (251, 201, 17), (252, 203, 8), (254, 202, 7), (252, 195, 0), (252, 192, 0), (253, 195, 0), (251, 177, 21), (238, 125, 55), (240, 117, 48), (241, 115, 8), (243, 109, 1), (241, 107, 1), (243, 106, 0), (242, 105, 0), (242, 105, 0), (242, 104, 1), (242, 104, 1), (244, 106, 2), (244, 106, 2), (243, 106, 1), (242, 105, 1), (242, 105, 1), (242, 105, 1), (243, 105, 1), (243, 104, 1), (244, 106, 2), (244, 106, 2), (243, 105, 2), (243, 105, 1), (243, 105, 1), (241, 103, 0), (241, 103, 0), (241, 103, 0), (242, 103, 0), (243, 103, 0), (244, 102, 0), (243, 100, 0), (243, 100, 1), (243, 101, 0), (243, 100, 0), (243, 100, 0), (243, 100, 0), (243, 100, 0), (243, 101, 0), (244, 102, 0), (244, 102, 0), (243, 101, 0), (243, 101, 0), (243, 101, 0), (243, 101, 0), (243, 101, 0), (244, 100, 2), (244, 100, 2), (243, 100, 3), (243, 100, 2), (244, 100, 2), (244, 100, 2), (244, 100, 2), (244, 100, 0), (245, 100, 0), (245, 99, 1), (245, 99, 1), (245, 99, 1), (245, 99, 1), (245, 99, 0), (246, 98, 2), (246, 97, 1), (246, 97, 2), (244, 96, 1), (244, 96, 1), (245, 94, 2), (245, 89, 2), (242, 82, 0), (240, 71, 3), (225, 28, 5), (208, 0, 0), (211, 1, 0), (212, 1, 1), (213, 2, 1), (214, 2, 0), (214, 2, 0), (213, 2, 0), (214, 2, 0), (215, 2, 0), (217, 2, 2), (217, 2, 2), (215, 1, 1), (215, 1, 1), (215, 1, 1), (215, 0, 1), (214, 1, 1), (214, 0, 0), (213, 0, 0), (212, 0, 0), (213, 0, 4), (212, 1, 10), (160, 124, 182), (164, 131, 187), (153, 120, 179), (129, 95, 161), (94, 60, 126), (49, 15, 77), (48, 17, 80), (58, 5, 73), (58, 0, 64), (69, 49, 90), (82, 56, 70), (62, 11, 16), (51, 11, 20), (41, 18, 27), (26, 9, 17), (26, 13, 31), (39, 19, 45), (37, 18, 42), (36, 15, 36), (36, 26, 48), (26, 109, 190), (0, 106, 209), (0, 90, 200), (2, 87, 201), (1, 81, 194), (1, 78, 191), (1, 75, 189), (0, 70, 186), (0, 66, 184), (0, 62, 183), (0, 62, 182), (1, 63, 178), (1, 63, 174), (1, 63, 172), (0, 64, 172), (0, 65, 175), (1, 66, 177), (2, 72, 180), (0, 78, 180), (0, 90, 200), (25, 91, 184), (30, 21, 36), (43, 20, 3), (66, 27, 5), (112, 50, 17), (215, 150, 27), (235, 171, 1), (236, 171, 2), (237, 171, 3), (236, 171, 1), (236, 171, 0), (237, 169, 0), (240, 168, 0), (241, 168, 0), (243, 167, 0), (244, 167, 0), (245, 166, 0), (246, 167, 0), (248, 169, 1), (251, 170, 0), (254, 172, 0), (253, 176, 0), (255, 178, 1), (254, 179, 1), (252, 179, 1), (253, 181, 0), (254, 185, 2), (254, 182, 2), (253, 179, 1), (254, 179, 1), (254, 177, 9), (238, 136, 43), (238, 116, 52), (240, 114, 15), (242, 109, 1), (242, 106, 1), (244, 106, 0), (242, 105, 0), (242, 105, 0), (242, 104, 1), (242, 104, 1), (243, 105, 2), (243, 105, 2), (243, 104, 2), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (243, 105, 2), (243, 105, 2), (243, 105, 1), (241, 103, 0), (241, 103, 0), (241, 103, 0), (241, 103, 0), (241, 103, 0), (242, 103, 0), (243, 103, 0), (244, 101, 1), (243, 100, 1), (243, 100, 0), (243, 100, 0), (243, 100, 0), (243, 100, 0), (243, 99, 0), (243, 99, 0), (242, 100, 0), (244, 101, 0), (244, 101, 0), (242, 100, 0), (243, 100, 0), (243, 99, 0), (242, 99, 0), (242, 100, 1), (243, 99, 2), (243, 100, 2), (243, 100, 2), (243, 99, 2), (243, 98, 1), (243, 98, 1), (244, 98, 1), (243, 98, 0), (244, 98, 0), (244, 98, 2), (244, 98, 2), (244, 98, 2), (245, 98, 2), (246, 97, 2), (244, 96, 1), (244, 96, 2), (244, 95, 2), (243, 93, 0), (243, 92, 0), (243, 89, 0), (241, 83, 1), (236, 75, 0), (234, 58, 1), (217, 18, 3), (204, 0, 1), (207, 0, 0), (210, 1, 1), (210, 1, 1), (210, 1, 0), (209, 2, 0), (209, 2, 0), (209, 2, 0), (211, 2, 1), (212, 2, 2), (212, 2, 1), (210, 1, 0), (210, 1, 1), (210, 1, 0), (210, 1, 0), (210, 0, 0), (210, 0, 0), (208, 0, 0), (206, 0, 0), (209, 0, 1), (209, 1, 3), (220, 207, 238), (221, 208, 238), (225, 212, 240), (226, 210, 240), (214, 191, 227), (168, 139, 184), (87, 64, 113), (70, 44, 97), (84, 39, 98), (82, 46, 96), (63, 35, 64), (81, 39, 64), (126, 84, 111), (113, 75, 96), (91, 52, 72), (51, 27, 43), (32, 16, 35), (35, 19, 39), (35, 12, 28), (33, 57, 100), (11, 114, 208), (2, 91, 192), (0, 84, 190), (0, 81, 186), (0, 70, 179), (0, 56, 173), (0, 51, 165), (6, 54, 168), (9, 59, 170), (9, 61, 162), (8, 61, 159), (4, 57, 156), (0, 50, 153), (0, 43, 151), (0, 43, 156), (0, 49, 155), (1, 51, 157), (3, 57, 163), (3, 61, 166), (1, 68, 172), (5, 91, 196), (54, 60, 99), (88, 29, 0), (91, 30, 2), (89, 47, 19), (200, 144, 30), (234, 165, 0), (232, 165, 2), (232, 165, 3), (232, 166, 2), (233, 165, 0), (234, 163, 0), (237, 162, 1), (238, 161, 1), (239, 160, 1), (239, 160, 0), (240, 159, 1), (242, 160, 1), (245, 161, 0), (247, 163, 1), (247, 164, 0), (249, 165, 0), (250, 166, 1), (253, 165, 1), (254, 161, 0), (253, 161, 0), (253, 174, 2), (252, 175, 0), (251, 172, 0), (252, 172, 0), (255, 176, 2), (242, 150, 36), (237, 116, 52), (239, 113, 16), (241, 109, 0), (243, 106, 1), (244, 106, 1), (242, 106, 1), (242, 105, 0), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (241, 103, 0), (241, 103, 0), (241, 103, 0), (241, 103, 0), (241, 103, 0), (242, 103, 0), (243, 103, 0), (244, 101, 1), (243, 100, 1), (243, 101, 0), (243, 100, 0), (243, 100, 0), (243, 100, 0), (242, 99, 0), (242, 99, 1), (242, 99, 1), (243, 100, 0), (243, 100, 0), (242, 99, 1), (242, 99, 0), (242, 99, 0), (242, 99, 0), (243, 99, 1), (243, 98, 2), (242, 98, 1), (242, 98, 1), (243, 97, 0), (243, 96, 0), (244, 95, 0), (244, 96, 0), (243, 96, 0), (242, 96, 0), (242, 95, 1), (242, 95, 1), (242, 95, 1), (243, 95, 1), (244, 94, 1), (244, 94, 1), (243, 93, 1), (242, 92, 1), (241, 90, 1), (240, 87, 0), (239, 82, 0), (238, 76, 1), (234, 66, 0), (230, 47, 1), (210, 13, 5), (202, 0, 2), (206, 0, 1), (207, 1, 1), (206, 0, 1), (205, 1, 0), (204, 1, 0), (205, 1, 0), (205, 1, 0), (207, 1, 0), (207, 1, 1), (207, 1, 0), (206, 0, 0), (206, 0, 1), (207, 0, 0), (208, 1, 1), (208, 1, 1), (208, 1, 1), (207, 1, 1), (205, 1, 1), (205, 1, 0), (208, 1, 0), (201, 187, 224), (204, 190, 227), (206, 192, 229), (206, 192, 227), (207, 190, 227), (216, 193, 235), (203, 177, 222), (183, 154, 203), (192, 157, 209), (175, 139, 189), (128, 90, 139), (119, 82, 116), (140, 105, 126), (117, 83, 103), (90, 56, 73), (64, 44, 54), (34, 21, 32), (28, 12, 26), (34, 13, 28), (29, 79, 141), (3, 101, 200), (2, 83, 185), (0, 76, 184), (0, 65, 171), (11, 65, 167), (47, 97, 172), (78, 136, 183), (95, 159, 197), (82, 163, 193), (65, 165, 191), (49, 159, 183), (53, 143, 173), (66, 118, 162), (53, 90, 148), (28, 62, 142), (6, 38, 134), (0, 34, 139), (0, 43, 151), (3, 47, 155), (3, 52, 157), (0, 70, 177), (40, 76, 145), (90, 31, 2), (84, 29, 1), (62, 109, 121), (176, 157, 54), (227, 158, 0), (227, 159, 2), (228, 160, 0), (229, 161, 0), (230, 160, 0), (231, 159, 0), (234, 158, 1), (235, 158, 1), (235, 156, 0), (235, 155, 0), (236, 155, 0), (238, 154, 0), (241, 154, 0), (244, 157, 0), (244, 157, 0), (244, 156, 0), (244, 155, 0), (245, 151, 1), (244, 147, 3), (243, 144, 2), (249, 160, 2), (254, 173, 1), (252, 171, 0), (252, 171, 0), (255, 173, 0), (250, 162, 15), (237, 118, 56), (239, 109, 28), (240, 107, 3), (240, 106, 2), (241, 105, 1), (242, 106, 2), (242, 105, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (241, 103, 0), (241, 103, 0), (242, 104, 1), (242, 104, 1), (242, 104, 1), (244, 104, 1), (243, 104, 0), (243, 102, 0), (243, 100, 0), (243, 100, 0), (243, 100, 0), (243, 100, 0), (243, 100, 0), (243, 100, 1), (243, 100, 3), (243, 100, 3), (242, 98, 2), (242, 99, 1), (242, 99, 1), (242, 97, 0), (241, 97, 1), (241, 97, 0), (242, 96, 0), (243, 96, 0), (243, 97, 1), (243, 97, 1), (243, 95, 0), (243, 95, 0), (243, 95, 0), (243, 95, 0), (242, 94, 0), (243, 94, 0), (242, 93, 0), (242, 93, 0), (242, 93, 0), (242, 93, 0), (243, 93, 1), (243, 92, 1), (242, 91, 1), (241, 89, 1), (238, 86, 1), (236, 81, 0), (235, 75, 0), (235, 68, 1), (231, 55, 0), (228, 51, 10), (204, 24, 15), (196, 0, 1), (205, 1, 3), (204, 1, 0), (202, 1, 0), (201, 1, 0), (202, 1, 0), (204, 0, 1), (205, 0, 1), (205, 0, 0), (205, 1, 1), (204, 1, 1), (205, 0, 1), (205, 0, 1), (205, 0, 1), (206, 1, 2), (207, 1, 2), (208, 1, 0), (209, 1, 0), (207, 2, 1), (205, 2, 1), (207, 2, 0), (183, 166, 215), (187, 170, 219), (190, 173, 219), (189, 173, 217), (187, 170, 214), (186, 165, 211), (194, 171, 215), (195, 169, 211), (182, 154, 198), (174, 141, 190), (158, 119, 177), (126, 89, 132), (122, 94, 109), (125, 99, 105), (104, 76, 85), (70, 52, 57), (43, 30, 32), (31, 0, 4), (53, 7, 13), (25, 87, 154), (0, 91, 196), (0, 70, 172), (4, 69, 166), (50, 119, 178), (92, 179, 205), (97, 210, 220), (88, 215, 223), (73, 210, 221), (47, 205, 212), (19, 197, 206), (6, 190, 200), (14, 182, 195), (33, 170, 185), (40, 164, 180), (40, 152, 166), (38, 115, 150), (20, 65, 141), (0, 31, 131), (0, 34, 138), (4, 41, 145), (0, 47, 152), (33, 92, 160), (109, 71, 33), (73, 37, 21), (20, 140, 168), (146, 141, 59), (227, 151, 0), (220, 155, 1), (225, 156, 0), (227, 156, 0), (228, 155, 0), (229, 155, 0), (230, 155, 1), (231, 155, 1), (231, 153, 0), (232, 151, 0), (233, 150, 0), (235, 150, 0), (237, 150, 0), (239, 149, 0), (240, 149, 1), (238, 146, 0), (239, 144, 1), (239, 141, 2), (235, 136, 2), (233, 134, 1), (237, 140, 1), (252, 165, 4), (253, 172, 0), (254, 169, 0), (255, 169, 0), (254, 170, 2), (242, 136, 39), (234, 106, 43), (239, 106, 8), (239, 105, 0), (241, 104, 0), (242, 104, 0), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (242, 104, 1), (241, 103, 0), (241, 103, 0), (241, 103, 0), (241, 103, 0), (241, 103, 0), (242, 104, 1), (242, 104, 1), (243, 104, 1), (244, 104, 1), (243, 104, 0), (243, 102, 0), (243, 100, 0), (243, 100, 0), (243, 100, 0), (243, 100, 0), (243, 100, 2), (243, 100, 3), (243, 99, 2), (242, 98, 2), (241, 97, 2), (241, 97, 1), (241, 97, 0), (241, 98, 1), (241, 95, 0), (241, 93, 0), (240, 94, 0), (240, 95, 0), (241, 95, 1), (241, 95, 1), (242, 93, 0), (242, 93, 0), (242, 93, 0), (242, 93, 1), (242, 92, 0), (241, 92, 0), (240, 91, 0), (240, 91, 1), (240, 91, 0), (242, 91, 0), (242, 90, 0), (240, 88, 0), (239, 87, 1), (238, 84, 1), (235, 79, 0), (234, 74, 0), (233, 68, 1), (231, 61, 1), (223, 46, 0), (239, 70, 29), (207, 34, 23), (191, 0, 0), (201, 2, 3), (199, 2, 1), (198, 2, 0), (197, 2, 0), (199, 1, 0), (203, 2, 1), (203, 2, 1), (203, 1, 2), (205, 0, 2), (203, 2, 1), (203, 2, 1), (203, 2, 1), (202, 2, 1), (203, 2, 1), (204, 1, 1), (205, 0, 1), (205, 1, 0), (205, 1, 0), (204, 1, 1), (205, 0, 1), (165, 146, 203), (168, 150, 205), (170, 153, 205), (169, 152, 202), (171, 152, 200), (171, 151, 199), (173, 150, 198), (174, 149, 194), (172, 144, 189), (141, 110, 155), (125, 88, 136), (113, 74, 117), (95, 68, 85), (105, 85, 87), (105, 75, 83), (85, 56, 64), (43, 26, 25), (34, 1, 0), (46, 13, 19), (16, 86, 160), (0, 72, 171), (24, 93, 163), (82, 175, 207), (96, 214, 224), (63, 212, 219), (42, 204, 211), (38, 202, 211), (34, 201, 211), (22, 196, 206), (10, 194, 206), (3, 190, 204), (0, 185, 199), (0, 176, 192), (0, 171, 187), (0, 167, 182), (6, 159, 171), (24, 146, 164), (29, 99, 148), (9, 40, 130), (0, 32, 134), (1, 38, 141), (14, 66, 145), (72, 135, 142), (27, 141, 172), (1, 175, 230), (108, 146, 115), (219, 142, 0), (214, 150, 0), (220, 150, 0), (224, 151, 1), (224, 153, 0), (226, 153, 1), (228, 152, 1), (229, 150, 1), (230, 149, 1), (231, 148, 1), (231, 146, 1), (232, 146, 1), (233, 144, 0), (234, 143, 0), (235, 142, 1), (233, 139, 1), (233, 136, 0), (231, 134, 0), (228, 131, 0), (228, 130, 0), (228, 128, 0), (235, 139, 1), (247, 164, 3), (255, 169, 3), (255, 166, 3), (255, 169, 0), (251, 156, 15), (231, 112, 41), (235, 104, 13), (238, 104, 0), (238, 103, 1), (239, 102, 0), (241, 103, 1), (241, 103, 1), (241, 103, 1), (241, 103, 1), (241, 103, 1), (241, 103, 1), (241, 103, 2), (242, 104, 3), (242, 104, 2), (242, 104, 1), (242, 104, 1), (241, 103, 0), (241, 103, 0), (241, 103, 0), (241, 103, 0), (242, 104, 1), (242, 104, 1), (244, 104, 1), (244, 104, 1), (246, 103, 1), (245, 102, 0), (244, 101, 0), (243, 100, 0), (243, 100, 0), (243, 100, 0), (243, 100, 0), (242, 99, 1), (242, 99, 1), (241, 98, 0), (240, 97, 1), (241, 95, 1), (242, 96, 0), (241, 95, 0), (240, 95, 0), (241, 95, 0), (240, 94, 0), (239, 93, 0), (239, 93, 0), (240, 92, 1), (241, 92, 0), (241, 92, 0), (240, 91, 0), (240, 91, 0), (240, 90, 1), (239, 90, 1), (239, 89, 0), (240, 88, 0), (240, 89, 2), (240, 88, 0), (240, 88, 0), (240, 88, 1), (239, 86, 2), (238, 83, 2), (235, 79, 1), (233, 74, 1), (233, 69, 2), (230, 63, 1), (225, 55, 0), (226, 49, 3), (246, 72, 29), (205, 27, 12), (189, 0, 1), (196, 0, 2), (194, 0, 0), (195, 0, 1), (197, 1, 1), (197, 0, 1), (201, 0, 1), (202, 1, 0), (203, 1, 1), (204, 1, 2), (204, 1, 1), (202, 1, 0), (201, 1, 0), (202, 1, 0), (204, 1, 1), (204, 1, 1), (204, 1, 1), (205, 0, 1), (206, 0, 1), (206, 0, 1), (205, 0, 1), (145, 127, 185), (149, 130, 189), (149, 132, 188), (150, 132, 185), (152, 131, 186), (153, 130, 185), (155, 128, 180), (153, 125, 174), (152, 122, 170), (137, 107, 145), (97, 67, 89), (97, 65, 91), (79, 53, 75), (71, 48, 63), (84, 54, 72), (85, 55, 73), (62, 37, 50), (38, 12, 22), (22, 12, 30), (6, 70, 153), (33, 116, 179), (87, 197, 214), (63, 209, 221), (22, 194, 203), (4, 188, 198), (0, 183, 195), (0, 180, 191), (0, 180, 190), (1, 180, 192), (2, 181, 196), (2, 184, 199), (3, 185, 199), (4, 177, 193), (2, 170, 187), (2, 168, 185), (0, 162, 177), (1, 155, 167), (13, 156, 166), (25, 121, 151), (9, 46, 136), (0, 29, 144), (0, 44, 139), (50, 174, 229), (8, 199, 255), (0, 185, 255), (53, 154, 176), (194, 133, 6), (214, 143, 0), (213, 146, 1), (219, 147, 1), (223, 150, 0), (225, 151, 1), (227, 149, 0), (227, 147, 1), (227, 145, 2), (229, 144, 2), (229, 143, 1), (229, 141, 1), (228, 140, 0), (230, 138, 0), (229, 136, 1), (229, 134, 1), (228, 131, 0), (226, 128, 1), (224, 126, 0), (223, 124, 0), (225, 124, 0), (230, 125, 1), (235, 134, 2), (242, 149, 2), (245, 152, 3), (246, 153, 3), (248, 150, 5), (233, 123, 31), (228, 102, 38), (235, 102, 4), (238, 100, 0), (238, 100, 0), (240, 102, 0), (240, 102, 0), (240, 102, 0), (240, 102, 0), (240, 102, 0), (240, 102, 0), (240, 102, 1), (241, 104, 3), (241, 103, 2), (241, 103, 0), (241, 103, 0), (241, 103, 0), (241, 103, 1), (241, 103, 1), (241, 103, 0), (242, 104, 1), (242, 104, 1), (244, 104, 1), (245, 103, 1), (246, 103, 1), (245, 102, 0), (244, 101, 0), (243, 100, 0), (243, 100, 0), (242, 99, 0), (242, 99, 0), (242, 100, 0), (243, 99, 2), (241, 97, 1), (241, 95, 2), (241, 95, 1), (241, 96, 0), (240, 94, 0), (240, 94, 0), (240, 94, 0), (239, 93, 0), (238, 92, 0), (238, 91, 1), (239, 92, 2), (239, 91, 1), (238, 89, 0), (238, 89, 0), (238, 88, 1), (238, 88, 1), (239, 88, 1), (240, 87, 1), (240, 87, 2), (239, 86, 1), (237, 84, 0), (237, 84, 0), (237, 84, 1), (237, 83, 2), (236, 79, 2), (233, 74, 2), (231, 69, 1), (229, 63, 2), (226, 58, 1), (222, 51, 1), (234, 61, 19), (236, 51, 13), (209, 14, 4), (187, 0, 1), (190, 1, 3), (190, 0, 1), (192, 1, 4), (195, 1, 3), (197, 1, 1), (199, 0, 1), (201, 2, 0), (201, 1, 0), (201, 1, 0), (201, 1, 0), (201, 0, 0), (200, 0, 0), (200, 0, 0), (201, 1, 0), (201, 1, 0), (202, 1, 0), (203, 0, 0), (202, 1, 0), (203, 0, 0), (203, 1, 0), (129, 110, 169), (132, 114, 174), (133, 114, 172), (134, 114, 169), (135, 112, 169), (138, 111, 167), (139, 108, 164), (136, 104, 156), (132, 99, 149), (133, 102, 138), (99, 72, 83), (82, 56, 73), (70, 43, 74), (114, 85, 124), (157, 123, 165), (165, 122, 166), (148, 108, 150), (126, 89, 128), (71, 52, 82), (48, 112, 153), (77, 205, 225), (30, 197, 205), (2, 181, 195), (0, 176, 186), (0, 170, 183), (0, 165, 182), (1, 162, 180), (1, 160, 176), (1, 160, 176), (1, 162, 180), (2, 166, 183), (3, 169, 187), (2, 170, 189), (3, 172, 189), (4, 171, 187), (2, 164, 181), (0, 157, 173), (1, 152, 167), (0, 150, 160), (1, 113, 143), (0, 46, 133), (14, 57, 151), (160, 196, 223), (140, 216, 238), (52, 178, 225), (46, 169, 205), (158, 132, 58), (207, 128, 0), (205, 138, 0), (216, 144, 0), (219, 148, 2), (223, 149, 2), (224, 147, 1), (224, 146, 0), (225, 143, 1), (224, 141, 1), (223, 139, 0), (224, 136, 0), (225, 135, 0), (225, 133, 0), (224, 131, 0), (222, 128, 0), (223, 126, 0), (223, 124, 2), (220, 121, 1), (219, 118, 1), (221, 119, 1), (226, 120, 3), (226, 123, 3), (228, 131, 2), (228, 131, 2), (231, 131, 2), (234, 131, 0), (233, 129, 10), (226, 110, 36), (233, 101, 13), (239, 100, 0), (239, 100, 2), (240, 101, 1), (240, 102, 1), (240, 102, 1), (240, 102, 1), (240, 102, 1), (240, 102, 1), (240, 102, 1), (241, 102, 2), (241, 103, 1), (241, 103, 0), (241, 103, 0), (241, 103, 1), (241, 103, 2), (241, 103, 2), (241, 103, 1), (242, 104, 1), (243, 104, 1), (245, 104, 1), (246, 103, 1), (246, 103, 1), (245, 102, 0), (244, 101, 0), (243, 100, 0), (243, 100, 0), (242, 99, 0), (242, 99, 1), (243, 100, 2), (243, 99, 3), (241, 97, 2), (242, 96, 2), (242, 95, 1), (240, 96, 1), (240, 95, 0), (240, 94, 0), (240, 93, 0), (238, 91, 0), (237, 90, 0), (238, 89, 1), (238, 90, 2), (238, 90, 1), (238, 88, 1), (238, 88, 1), (239, 88, 2), (239, 87, 3), (240, 87, 2), (240, 86, 2), (238, 86, 3), (237, 84, 2), (234, 82, 0), (234, 82, 1), (235, 81, 2), (234, 80, 2), (233, 75, 2), (230, 70, 2), (228, 64, 1), (226, 57, 0), (230, 52, 0), (209, 49, 8), (214, 58, 30), (222, 20, 7), (208, 0, 0), (189, 2, 0), (187, 1, 2), (187, 0, 2), (189, 0, 3), (192, 1, 1), (194, 2, 1), (197, 1, 1), (198, 2, 0), (199, 2, 0), (199, 1, 1), (199, 1, 1), (199, 0, 0), (198, 0, 0), (198, 1, 0), (199, 2, 1), (199, 2, 1), (201, 1, 0), (201, 1, 0), (200, 2, 0), (201, 1, 0), (201, 1, 0), (112, 93, 152), (115, 95, 155), (117, 94, 153), (118, 95, 151), (121, 95, 151), (123, 95, 149), (124, 95, 148), (124, 96, 139), (122, 93, 128), (122, 94, 119), (100, 75, 82), (66, 40, 57), (108, 81, 118), (167, 137, 188), (168, 135, 183), (161, 156, 190), (158, 198, 216), (143, 217, 224), (115, 198, 206), (60, 189, 198), (15, 188, 194), (3, 173, 186), (1, 164, 180), (0, 159, 171), (0, 154, 166), (0, 150, 166), (0, 149, 165), (1, 147, 163), (2, 147, 164), (1, 149, 168), (0, 150, 170), (1, 153, 173), (1, 157, 177), (2, 162, 180), (4, 165, 183), (3, 164, 183), (0, 157, 174), (0, 140, 163), (18, 151, 168), (103, 183, 189), (172, 206, 221), (208, 229, 235), (229, 247, 250), (238, 250, 255), (237, 245, 251), (223, 244, 250), (214, 228, 222), (217, 195, 152), (208, 158, 65), (206, 133, 2), (215, 138, 0), (220, 146, 1), (220, 145, 1), (222, 145, 1), (221, 141, 0), (220, 138, 0), (219, 136, 0), (220, 133, 0), (221, 131, 0), (219, 129, 1), (218, 127, 1), (216, 124, 0), (217, 122, 0), (218, 120, 1), (216, 117, 0), (214, 114, 2), (217, 113, 2), (216, 112, 4), (218, 119, 3), (224, 128, 2), (226, 129, 3), (229, 130, 3), (230, 130, 0), (231, 132, 3), (226, 119, 21), (228, 101, 27), (234, 97, 6), (236, 98, 1), (239, 101, 2), (239, 101, 2), (239, 100, 2), (239, 100, 2), (239, 100, 2), (240, 101, 2), (240, 101, 2), (240, 101, 2), (240, 102, 1), (240, 102, 0), (240, 102, 0), (241, 103, 2), (241, 103, 2), (241, 103, 2), (241, 103, 2), (242, 103, 2), (244, 103, 1), (246, 103, 1), (246, 103, 1), (246, 103, 1), (245, 103, 0), (243, 101, 0), (242, 99, 0), (242, 99, 0), (243, 100, 0), (243, 100, 2), (243, 99, 2), (241, 97, 2), (241, 97, 2), (242, 97, 2), (243, 96, 2), (241, 95, 1), (240, 94, 0), (240, 94, 0), (239, 93, 0), (238, 91, 0), (238, 89, 0), (238, 88, 0), (237, 88, 0), (237, 88, 1), (238, 86, 2), (238, 85, 1), (238, 85, 1), (237, 84, 2), (237, 84, 2), (237, 84, 2), (236, 82, 2), (235, 82, 2), (234, 81, 2), (233, 80, 2), (232, 78, 3), (230, 75, 3), (229, 70, 2), (227, 64, 0), (224, 57, 0), (227, 53, 0), (216, 54, 4), (121, 46, 12), (193, 41, 18), (213, 5, 0), (205, 0, 2), (191, 2, 0), (187, 0, 1), (186, 0, 2), (187, 0, 2), (189, 0, 0), (192, 1, 0), (195, 2, 1), (196, 1, 0), (198, 1, 1), (199, 1, 2), (199, 1, 2), (198, 0, 1), (197, 1, 1), (196, 1, 1), (197, 1, 1), (199, 1, 1), (200, 1, 0), (200, 1, 0), (200, 1, 1), (200, 1, 0), (200, 1, 0), (99, 81, 128), (102, 82, 132), (103, 80, 131), (104, 80, 130), (109, 84, 133), (113, 87, 129), (114, 88, 126), (113, 89, 118), (110, 91, 106), (113, 94, 98), (84, 61, 66), (56, 29, 49), (118, 87, 125), (133, 100, 145), (136, 140, 169), (126, 231, 232), (74, 240, 234), (55, 226, 222), (53, 204, 210), (12, 181, 186), (0, 166, 175), (2, 157, 167), (0, 147, 159), (0, 142, 153), (1, 140, 150), (1, 136, 150), (1, 134, 148), (1, 134, 147), (2, 136, 152), (2, 136, 155), (2, 138, 158), (1, 142, 160), (0, 145, 162), (1, 149, 167), (1, 154, 173), (0, 153, 176), (3, 148, 168), (97, 188, 198), (202, 237, 244), (245, 251, 255), (239, 255, 255), (233, 251, 255), (228, 246, 253), (227, 246, 252), (229, 245, 254), (232, 246, 255), (228, 250, 255), (228, 252, 255), (233, 243, 250), (219, 207, 176), (205, 152, 53), (210, 134, 0), (218, 142, 0), (218, 142, 1), (217, 140, 1), (217, 136, 1), (215, 134, 1), (215, 131, 0), (215, 128, 0), (213, 125, 0), (212, 124, 0), (211, 121, 0), (211, 119, 0), (210, 117, 0), (207, 114, 0), (206, 112, 0), (209, 113, 3), (174, 86, 9), (199, 111, 6), (221, 126, 2), (219, 125, 2), (223, 128, 2), (225, 129, 2), (226, 128, 3), (224, 123, 6), (221, 110, 24), (228, 98, 22), (234, 96, 3), (237, 98, 2), (238, 99, 3), (238, 99, 2), (239, 100, 0), (239, 100, 1), (240, 101, 2), (240, 101, 2), (240, 101, 2), (240, 102, 1), (240, 102, 0), (240, 102, 0), (240, 102, 0), (240, 102, 0), (240, 102, 0), (240, 102, 0), (241, 101, 0), (243, 102, 0), (244, 102, 0), (244, 102, 0), (244, 102, 0), (243, 101, 0), (243, 99, 0), (242, 99, 0), (242, 99, 0), (242, 99, 2), (242, 99, 1), (242, 99, 0), (241, 97, 1), (242, 98, 0), (242, 97, 0), (241, 95, 0), (240, 94, 0), (240, 94, 0), (240, 93, 0), (239, 92, 1), (237, 90, 2), (236, 88, 1), (236, 87, 0), (236, 86, 0), (236, 86, 1), (238, 86, 3), (238, 85, 3), (235, 82, 1), (234, 80, 1), (234, 80, 1), (233, 80, 1), (233, 79, 1), (232, 78, 2), (232, 76, 1), (230, 75, 1), (228, 72, 2), (226, 69, 2), (225, 63, 0), (224, 57, 0), (222, 52, 0), (226, 52, 6), (131, 41, 10), (50, 31, 11), (168, 24, 10), (203, 0, 0), (195, 0, 0), (186, 0, 0), (183, 0, 0), (186, 1, 0), (185, 1, 1), (187, 1, 0), (191, 1, 0), (193, 1, 0), (194, 0, 0), (195, 1, 0), (195, 2, 1), (195, 2, 1), (195, 2, 1), (195, 2, 1), (195, 2, 1), (195, 2, 1), (195, 1, 1), (197, 1, 1), (197, 1, 1), (197, 1, 1), (198, 2, 0), (198, 2, 0), (88, 70, 106), (91, 70, 107), (92, 70, 107), (95, 71, 110), (98, 73, 114), (102, 79, 112), (101, 82, 104), (103, 85, 100), (103, 79, 86), (104, 86, 82), (104, 98, 96), (94, 100, 112), (108, 113, 127), (90, 89, 103), (88, 186, 188), (25, 223, 217), (0, 206, 204), (20, 194, 201), (19, 177, 188), (1, 159, 169), (1, 147, 158), (0, 138, 148), (0, 131, 143), (1, 126, 140), (1, 125, 138), (2, 122, 138), (2, 122, 137), (2, 123, 137), (3, 123, 140), (3, 125, 144), (1, 129, 146), (1, 131, 150), (1, 134, 153), (1, 137, 156), (0, 136, 160), (17, 146, 168), (153, 214, 229), (238, 251, 255), (229, 243, 255), (214, 238, 254), (211, 236, 254), (211, 235, 253), (212, 235, 251), (208, 234, 250), (204, 233, 251), (209, 233, 251), (211, 234, 253), (213, 235, 254), (218, 240, 254), (226, 249, 255), (228, 235, 237), (205, 164, 83), (210, 128, 0), (217, 138, 3), (214, 135, 2), (211, 131, 1), (209, 128, 1), (211, 126, 1), (208, 123, 0), (207, 120, 0), (207, 120, 1), (206, 117, 0), (206, 115, 0), (204, 113, 0), (203, 110, 0), (207, 110, 4), (174, 88, 10), (118, 51, 3), (180, 100, 8), (214, 124, 3), (215, 124, 4), (218, 124, 2), (219, 125, 0), (221, 124, 1), (218, 121, 0), (216, 114, 7), (225, 98, 30), (233, 93, 15), (234, 95, 1), (236, 96, 2), (237, 97, 2), (237, 98, 1), (239, 100, 3), (239, 100, 1), (239, 100, 1), (240, 101, 2), (240, 102, 1), (240, 102, 0), (240, 102, 0), (241, 102, 0), (242, 101, 0), (242, 101, 2), (242, 102, 3), (243, 102, 2), (243, 102, 1), (243, 102, 0), (243, 102, 1), (243, 102, 2), (243, 102, 2), (243, 101, 1), (242, 99, 1), (242, 99, 1), (242, 99, 1), (242, 98, 1), (241, 97, 0), (242, 97, 0), (243, 97, 0), (242, 95, 0), (241, 95, 1), (240, 94, 0), (239, 93, 0), (238, 92, 1), (238, 90, 1), (238, 88, 2), (236, 87, 1), (234, 85, 0), (234, 84, 0), (234, 83, 0), (235, 82, 1), (235, 82, 2), (234, 81, 2), (233, 79, 1), (232, 78, 0), (231, 77, 0), (230, 75, 0), (230, 73, 1), (228, 70, 0), (226, 68, 0), (225, 66, 2), (222, 63, 1), (222, 57, 1), (220, 52, 0), (224, 53, 4), (147, 38, 10), (48, 18, 3), (66, 26, 7), (156, 36, 19), (214, 28, 26), (219, 43, 39), (227, 56, 51), (195, 23, 19), (178, 0, 0), (185, 1, 1), (187, 0, 1), (191, 1, 2), (193, 0, 2), (196, 1, 3), (195, 0, 1), (194, 0, 0), (194, 0, 0), (195, 2, 1), (195, 2, 1), (196, 1, 1), (195, 0, 0), (194, 0, 0), (195, 0, 0), (195, 0, 0), (195, 0, 0), (196, 1, 0), (196, 1, 0), (80, 62, 87), (82, 62, 88), (83, 62, 88), (87, 65, 89), (89, 67, 90), (93, 72, 90), (95, 77, 88), (94, 75, 73), (108, 109, 103), (151, 199, 188), (161, 245, 238), (153, 253, 250), (145, 243, 239), (129, 223, 224), (63, 214, 211), (0, 188, 184), (5, 186, 188), (21, 180, 186), (2, 157, 163), (0, 143, 152), (1, 130, 141), (0, 121, 132), (1, 116, 127), (2, 112, 126), (2, 110, 124), (2, 110, 124), (2, 110, 124), (1, 110, 124), (0, 112, 127), (1, 115, 131), (1, 118, 135), (2, 121, 138), (2, 124, 142), (0, 125, 143), (11, 132, 150), (157, 220, 227), (228, 246, 254), (203, 233, 251), (195, 229, 250), (193, 227, 249), (187, 225, 249), (186, 222, 246), (183, 221, 248), (175, 217, 248), (174, 217, 247), (178, 220, 248), (185, 222, 249), (192, 225, 252), (199, 229, 253), (206, 232, 250), (214, 239, 255), (221, 235, 247), (207, 156, 86), (208, 120, 0), (207, 131, 2), (204, 126, 1), (203, 123, 0), (203, 121, 1), (202, 118, 1), (201, 115, 1), (201, 113, 2), (199, 111, 0), (199, 109, 0), (199, 108, 0), (199, 109, 6), (167, 88, 8), (122, 54, 6), (114, 52, 1), (173, 91, 6), (203, 119, 3), (204, 119, 2), (208, 119, 2), (211, 120, 0), (211, 117, 0), (210, 113, 1), (207, 110, 1), (209, 103, 19), (218, 96, 33), (227, 92, 14), (235, 94, 0), (235, 95, 1), (235, 95, 1), (237, 97, 2), (237, 98, 1), (238, 99, 1), (239, 100, 2), (239, 100, 1), (239, 100, 1), (240, 100, 1), (242, 100, 3), (242, 101, 2), (242, 101, 3), (243, 102, 4), (243, 102, 4), (242, 101, 2), (242, 101, 0), (242, 101, 0), (242, 101, 3), (242, 102, 3), (242, 100, 1), (242, 99, 0), (242, 99, 0), (242, 99, 1), (242, 98, 1), (242, 96, 1), (243, 97, 2), (241, 95, 0), (240, 94, 0), (240, 93, 2), (239, 92, 1), (238, 91, 1), (237, 89, 1), (236, 88, 1), (235, 86, 0), (235, 85, 0), (233, 83, 0), (233, 82, 0), (231, 81, 0), (233, 79, 1), (233, 79, 1), (233, 79, 1), (231, 78, 0), (229, 76, 0), (228, 74, 0), (228, 71, 1), (228, 69, 1), (227, 65, 0), (225, 63, 0), (224, 62, 1), (220, 57, 0), (218, 53, 0), (222, 50, 4), (180, 44, 10), (108, 36, 13), (153, 46, 32), (193, 59, 44), (210, 68, 47), (223, 74, 60), (232, 83, 72), (239, 92, 80), (226, 75, 65), (181, 8, 8), (182, 0, 0), (186, 1, 2), (188, 2, 3), (191, 1, 1), (193, 1, 3), (195, 0, 1), (195, 0, 0), (194, 0, 0), (195, 2, 1), (195, 2, 1), (195, 1, 1), (195, 0, 0), (195, 0, 0), (195, 0, 0), (195, 0, 0), (195, 0, 0), (195, 0, 0), (195, 0, 0), (77, 62, 70), (76, 64, 72), (75, 61, 72), (81, 63, 74), (86, 66, 74), (91, 70, 71), (99, 70, 58), (103, 109, 87), (132, 229, 224), (101, 249, 247), (67, 239, 238), (53, 235, 233), (52, 233, 237), (58, 240, 243), (75, 240, 246), (32, 200, 206), (10, 168, 176), (12, 165, 172), (0, 142, 149), (3, 125, 135), (3, 115, 127), (3, 108, 119), (2, 105, 116), (1, 103, 114), (1, 101, 113), (2, 101, 113), (2, 101, 113), (1, 102, 114), (0, 104, 117), (0, 106, 121), (1, 109, 125), (1, 113, 129), (1, 116, 133), (0, 111, 128), (120, 189, 208), (212, 239, 255), (191, 225, 246), (179, 217, 247), (170, 212, 242), (165, 209, 238), (161, 208, 241), (156, 207, 244), (144, 200, 241), (144, 200, 242), (146, 202, 241), (152, 206, 243), (161, 208, 246), (169, 211, 248), (178, 215, 248), (186, 221, 249), (196, 223, 250), (204, 231, 255), (208, 226, 234), (187, 131, 43), (197, 116, 0), (201, 121, 1), (198, 119, 3), (197, 115, 2), (197, 113, 2), (196, 110, 3), (193, 108, 1), (194, 107, 0), (196, 106, 1), (183, 98, 9), (125, 69, 23), (69, 35, 27), (107, 54, 9), (163, 81, 3), (183, 91, 3), (182, 98, 1), (190, 107, 2), (196, 111, 2), (198, 111, 1), (202, 108, 1), (199, 104, 4), (198, 100, 3), (213, 113, 2), (226, 120, 20), (220, 94, 29), (229, 89, 7), (231, 91, 0), (231, 92, 0), (234, 94, 2), (235, 95, 2), (235, 96, 2), (237, 97, 1), (237, 98, 0), (238, 99, 1), (240, 99, 3), (240, 99, 3), (239, 99, 3), (239, 100, 2), (241, 101, 2), (241, 101, 2), (242, 101, 2), (242, 101, 2), (242, 101, 2), (242, 100, 2), (242, 100, 1), (243, 100, 0), (243, 100, 0), (243, 100, 1), (242, 99, 2), (242, 99, 1), (242, 97, 1), (242, 96, 3), (240, 95, 1), (238, 93, 0), (239, 91, 2), (238, 90, 1), (237, 89, 2), (236, 88, 1), (235, 86, 0), (234, 85, 0), (234, 83, 1), (234, 81, 1), (232, 79, 0), (229, 78, 1), (230, 76, 1), (229, 75, 1), (229, 74, 1), (228, 74, 1), (227, 73, 0), (225, 71, 0), (225, 68, 1), (224, 65, 1), (224, 62, 2), (223, 59, 1), (220, 56, 0), (218, 53, 0), (217, 49, 2), (204, 37, 5), (180, 24, 7), (198, 32, 10), (211, 38, 14), (210, 41, 21), (207, 47, 31), (206, 52, 38), (210, 57, 45), (212, 58, 49), (217, 65, 57), (203, 41, 38), (178, 2, 2), (181, 1, 1), (184, 3, 2), (188, 1, 1), (190, 2, 1), (193, 1, 1), (195, 0, 1), (194, 0, 1), (194, 2, 1), (194, 2, 1), (196, 2, 0), (197, 0, 0), (197, 1, 0), (197, 0, 2), (193, 0, 2), (193, 1, 2), (195, 0, 1), (195, 0, 1), (80, 64, 63), (90, 70, 63), (87, 63, 52), (79, 58, 44), (80, 62, 45), (93, 73, 42), (100, 83, 37), (93, 179, 162), (29, 224, 227), (0, 209, 217), (0, 214, 220), (0, 216, 220), (0, 216, 222), (0, 216, 219), (8, 214, 215), (15, 218, 221), (8, 176, 185), (5, 142, 153), (2, 125, 136), (3, 112, 121), (2, 103, 113), (1, 100, 109), (0, 97, 107), (0, 94, 105), (0, 93, 104), (1, 93, 105), (1, 94, 105), (0, 96, 107), (0, 98, 111), (0, 100, 114), (0, 102, 118), (1, 105, 122), (0, 100, 118), (52, 136, 157), (192, 228, 251), (182, 212, 237), (165, 204, 232), (150, 200, 235), (139, 195, 235), (133, 191, 237), (130, 189, 238), (120, 184, 236), (112, 185, 234), (115, 186, 235), (117, 187, 237), (127, 190, 238), (138, 195, 241), (147, 195, 240), (158, 199, 240), (168, 205, 244), (179, 211, 246), (186, 213, 247), (195, 225, 255), (195, 180, 167), (174, 99, 5), (193, 109, 0), (194, 114, 2), (194, 113, 2), (192, 109, 0), (186, 105, 0), (180, 104, 2), (169, 98, 11), (136, 76, 21), (82, 49, 36), (47, 33, 51), (59, 32, 43), (138, 71, 19), (174, 88, 4), (172, 85, 1), (171, 86, 1), (172, 90, 2), (177, 94, 3), (182, 97, 3), (184, 97, 3), (183, 93, 2), (188, 90, 1), (209, 109, 2), (225, 124, 5), (218, 108, 21), (218, 86, 28), (227, 84, 8), (227, 88, 0), (230, 90, 1), (232, 91, 1), (233, 93, 1), (234, 95, 1), (235, 95, 0), (235, 96, 1), (236, 97, 1), (237, 97, 2), (237, 97, 1), (237, 97, 1), (238, 99, 2), (238, 101, 1), (240, 100, 1), (241, 99, 2), (241, 100, 1), (241, 99, 1), (243, 100, 0), (244, 101, 1), (244, 101, 2), (244, 101, 2), (243, 100, 2), (243, 100, 2), (242, 99, 1), (241, 97, 2), (239, 95, 0), (238, 92, 1), (238, 90, 2), (237, 88, 1), (237, 87, 1), (236, 87, 0), (234, 84, 0), (233, 81, 0), (231, 80, 1), (232, 78, 1), (230, 76, 0), (227, 74, 0), (227, 73, 0), (226, 71, 0), (224, 69, 0), (224, 69, 0), (224, 70, 0), (224, 67, 0), (222, 64, 1), (220, 62, 1), (220, 58, 2), (220, 56, 1), (219, 51, 2), (218, 48, 4), (201, 27, 5), (180, 3, 1), (183, 0, 1), (186, 3, 2), (185, 11, 0), (189, 16, 4), (193, 23, 12), (194, 27, 14), (194, 29, 17), (196, 28, 19), (193, 23, 16), (189, 24, 16), (176, 5, 4), (174, 0, 1), (181, 1, 1), (185, 1, 1), (189, 2, 1), (191, 1, 1), (193, 1, 2), (194, 0, 2), (192, 1, 0), (193, 2, 1), (197, 2, 0), (200, 1, 0), (199, 2, 1), (198, 1, 4), (191, 1, 3), (191, 2, 4), (194, 2, 3), (194, 1, 3), (78, 62, 47), (84, 69, 38), (97, 86, 60), (118, 122, 114), (150, 159, 155), (170, 182, 170), (175, 194, 182), (151, 224, 233), (105, 220, 230), (65, 212, 216), (26, 198, 216), (0, 193, 207), (0, 193, 203), (0, 196, 205), (0, 193, 203), (2, 193, 205), (3, 169, 179), (4, 129, 139), (4, 113, 123), (3, 103, 111), (1, 94, 103), (0, 92, 99), (0, 90, 98), (1, 87, 97), (1, 86, 96), (1, 87, 97), (1, 88, 97), (1, 89, 99), (1, 92, 103), (1, 91, 104), (1, 93, 107), (1, 97, 111), (0, 90, 105), (120, 179, 203), (181, 216, 245), (150, 196, 224), (126, 186, 228), (105, 179, 231), (100, 175, 230), (97, 171, 229), (93, 169, 229), (84, 165, 230), (84, 168, 232), (88, 170, 231), (95, 170, 233), (104, 174, 233), (116, 180, 233), (126, 182, 233), (136, 186, 235), (147, 191, 237), (158, 196, 238), (167, 199, 240), (175, 206, 248), (189, 211, 243), (116, 99, 83), (104, 66, 13), (125, 82, 15), (130, 86, 11), (128, 82, 10), (119, 70, 5), (99, 57, 25), (62, 45, 56), (49, 36, 68), (50, 38, 69), (58, 38, 71), (105, 61, 36), (156, 83, 9), (160, 80, 0), (163, 84, 1), (164, 85, 2), (161, 83, 1), (159, 82, 0), (165, 84, 1), (170, 85, 0), (175, 87, 0), (183, 90, 0), (199, 102, 0), (211, 112, 1), (210, 110, 4), (199, 92, 16), (211, 83, 15), (221, 84, 2), (225, 87, 0), (227, 88, 0), (230, 90, 0), (232, 92, 0), (232, 92, 1), (232, 93, 0), (233, 94, 0), (235, 96, 1), (234, 95, 1), (235, 96, 0), (237, 98, 1), (238, 99, 2), (238, 97, 2), (239, 97, 2), (239, 97, 0), (239, 98, 0), (238, 100, 1), (240, 101, 1), (243, 100, 2), (243, 100, 1), (242, 99, 1), (242, 98, 1), (241, 97, 0), (241, 95, 1), (237, 93, 1), (235, 93, 1), (235, 90, 2), (234, 88, 1), (233, 87, 1), (231, 85, 1), (230, 83, 1), (231, 80, 1), (229, 77, 0), (227, 75, 0), (227, 73, 0), (227, 72, 1), (225, 70, 1), (224, 69, 0), (221, 66, 0), (221, 66, 1), (221, 65, 2), (219, 63, 1), (219, 59, 1), (216, 57, 1), (215, 53, 0), (215, 51, 0), (214, 47, 7), (193, 25, 8), (169, 0, 1), (169, 0, 3), (172, 0, 3), (174, 1, 2), (174, 0, 1), (176, 1, 1), (177, 2, 0), (178, 2, 0), (175, 4, 0), (173, 3, 0), (170, 0, 0), (168, 0, 0), (161, 1, 0), (157, 2, 0), (168, 1, 1), (182, 3, 1), (189, 1, 1), (189, 1, 1), (191, 2, 2), (192, 1, 2), (194, 0, 0), (194, 0, 0), (195, 1, 1), (198, 2, 2), (199, 2, 2), (197, 1, 1), (188, 1, 1), (189, 1, 3), (190, 2, 2), (191, 1, 2), (84, 76, 55), (147, 156, 145), (197, 218, 222), (216, 244, 255), (220, 249, 255), (216, 248, 255), (216, 245, 255), (217, 239, 255), (220, 239, 255), (212, 241, 255), (181, 233, 249), (117, 212, 233), (34, 185, 207), (0, 169, 188), (1, 168, 187), (2, 167, 188), (3, 150, 162), (0, 121, 129), (3, 104, 115), (2, 95, 105), (0, 89, 98), (0, 87, 94), (1, 85, 93), (1, 83, 92), (0, 81, 91), (0, 81, 92), (0, 82, 93), (1, 83, 94), (2, 84, 96), (1, 84, 97), (0, 86, 99), (0, 86, 100), (15, 98, 115), (139, 196, 222), (144, 192, 227), (114, 176, 223), (86, 166, 223), (65, 159, 225), (59, 156, 220), (59, 154, 218), (61, 151, 218), (52, 150, 220), (40, 148, 223), (50, 152, 224), (67, 153, 227), (79, 154, 224), (88, 158, 226), (98, 161, 226), (112, 166, 228), (122, 170, 231), (136, 175, 232), (150, 182, 234), (160, 189, 237), (176, 207, 249), (102, 131, 167), (16, 41, 55), (30, 49, 56), (34, 48, 55), (41, 44, 52), (52, 40, 39), (54, 39, 49), (44, 37, 71), (43, 41, 74), (57, 44, 78), (72, 44, 65), (132, 73, 12), (153, 77, 4), (158, 81, 3), (162, 85, 0), (162, 87, 0), (162, 87, 1), (163, 86, 1), (166, 86, 1), (174, 88, 1), (180, 91, 0), (186, 95, 0), (194, 100, 0), (200, 104, 1), (202, 103, 2), (192, 92, 0), (188, 82, 6), (209, 81, 10), (223, 81, 5), (226, 84, 0), (227, 86, 1), (230, 89, 2), (230, 89, 2), (231, 90, 1), (232, 92, 0), (233, 93, 1), (234, 94, 1), (234, 95, 1), (235, 96, 2), (236, 96, 1), (235, 96, 0), (235, 96, 1), (235, 96, 0), (235, 96, 0), (236, 97, 1), (238, 97, 1), (239, 97, 0), (239, 97, 0), (240, 96, 1), (239, 95, 0), (239, 95, 0), (238, 93, 1), (235, 90, 1), (234, 89, 1), (232, 87, 1), (231, 85, 0), (230, 85, 1), (229, 83, 1), (227, 80, 2), (227, 78, 2), (225, 75, 0), (224, 73, 1), (224, 72, 1), (224, 70, 1), (222, 68, 2), (219, 66, 2), (218, 64, 0), (218, 62, 1), (217, 61, 1), (216, 58, 1), (215, 55, 1), (213, 52, 2), (214, 49, 1), (208, 43, 4), (181, 18, 5), (161, 0, 0), (161, 2, 0), (162, 2, 1), (163, 2, 1), (166, 1, 0), (169, 1, 1), (169, 1, 1), (168, 1, 2), (167, 0, 3), (165, 0, 1), (162, 0, 0), (159, 0, 0), (156, 1, 0), (150, 1, 0), (144, 2, 0), (145, 1, 0), (156, 2, 2), (175, 2, 2), (187, 2, 2), (191, 3, 2), (193, 1, 2), (193, 1, 1), (193, 1, 1), (193, 1, 0), (195, 1, 0), (197, 1, 1), (198, 0, 2), (191, 2, 2), (190, 1, 1), (189, 1, 3), (188, 2, 1), (190, 205, 222), (217, 243, 255), (208, 241, 255), (199, 234, 255), (196, 231, 254), (193, 232, 255), (193, 231, 255), (193, 230, 254), (192, 229, 254), (194, 228, 254), (194, 230, 249), (198, 232, 253), (175, 228, 252), (79, 190, 213), (0, 149, 170), (0, 149, 170), (6, 138, 152), (0, 113, 121), (2, 97, 107), (2, 90, 98), (0, 84, 92), (0, 82, 88), (0, 80, 87), (0, 77, 87), (0, 75, 84), (0, 77, 84), (0, 78, 86), (0, 79, 89), (2, 80, 91), (1, 80, 91), (1, 80, 91), (0, 75, 84), (33, 105, 128), (125, 184, 224), (107, 166, 222), (80, 158, 218), (53, 150, 217), (27, 143, 217), (13, 141, 213), (15, 139, 212), (21, 131, 206), (37, 135, 212), (29, 133, 215), (17, 133, 214), (27, 135, 217), (50, 135, 218), (68, 137, 222), (79, 142, 224), (95, 147, 225), (109, 152, 229), (120, 158, 230), (131, 164, 230), (139, 172, 230), (158, 187, 242), (126, 160, 203), (10, 60, 79), (17, 60, 78), (26, 58, 77), (37, 53, 71), (50, 48, 60), (57, 45, 47), (50, 42, 65), (49, 48, 81), (45, 42, 82), (80, 50, 38), (138, 77, 3), (146, 77, 4), (153, 82, 1), (158, 86, 0), (160, 87, 0), (163, 87, 0), (166, 87, 0), (170, 90, 0), (175, 92, 0), (180, 96, 0), (185, 97, 0), (190, 100, 0), (194, 102, 1), (193, 99, 1), (187, 90, 0), (183, 80, 2), (186, 76, 8), (199, 75, 14), (216, 76, 6), (224, 81, 1), (225, 84, 1), (226, 85, 1), (228, 87, 1), (228, 88, 0), (230, 90, 1), (232, 92, 1), (232, 92, 1), (233, 93, 1), (233, 93, 0), (233, 94, 0), (233, 94, 1), (233, 94, 0), (233, 94, 0), (234, 95, 1), (235, 95, 1), (236, 94, 0), (236, 94, 1), (236, 94, 1), (233, 92, 0), (234, 92, 0), (235, 90, 1), (234, 88, 1), (232, 86, 1), (229, 84, 0), (228, 82, 0), (227, 81, 0), (226, 79, 2), (224, 76, 1), (224, 74, 0), (222, 72, 0), (221, 70, 1), (220, 67, 2), (219, 66, 1), (217, 63, 2), (215, 61, 2), (214, 59, 1), (213, 56, 0), (212, 55, 2), (210, 54, 2), (212, 51, 1), (212, 47, 3), (201, 34, 6), (173, 10, 3), (156, 0, 1), (156, 0, 0), (156, 1, 0), (157, 1, 0), (158, 1, 0), (159, 1, 0), (160, 1, 0), (160, 1, 0), (159, 1, 1), (156, 2, 1), (152, 2, 0), (150, 2, 0), (147, 2, 0), (145, 2, 1), (144, 1, 1), (142, 1, 1), (136, 1, 1), (134, 1, 2), (141, 1, 2), (154, 3, 2), (173, 3, 2), (186, 2, 0), (189, 2, 2), (192, 2, 1), (193, 2, 0), (193, 0, 1), (195, 0, 2), (200, 0, 4), (192, 2, 4), (188, 2, 3), (185, 1, 2), (185, 1, 0), (197, 234, 255), (190, 224, 246), (189, 224, 246), (184, 224, 248), (181, 223, 248), (178, 223, 249), (176, 221, 250), (176, 220, 249), (175, 219, 250), (171, 219, 249), (168, 218, 249), (168, 217, 247), (175, 218, 245), (174, 221, 254), (84, 185, 216), (2, 140, 162), (2, 133, 149), (0, 108, 116), (2, 93, 102), (2, 86, 93), (0, 81, 81), (0, 74, 76), (0, 70, 76), (0, 69, 79), (0, 70, 81), (0, 72, 79), (0, 71, 77), (0, 69, 77), (1, 72, 78), (1, 75, 83), (0, 76, 87), (0, 69, 76), (38, 110, 139), (94, 167, 224), (78, 146, 214), (57, 141, 205), (31, 137, 205), (6, 129, 203), (0, 128, 204), (0, 125, 202), (14, 124, 200), (35, 123, 206), (52, 121, 207), (43, 122, 205), (39, 122, 207), (47, 126, 210), (61, 127, 213), (75, 132, 216), (90, 135, 217), (102, 140, 220), (111, 146, 222), (118, 152, 223), (125, 158, 223), (141, 170, 234), (126, 162, 211), (7, 69, 84), (2, 62, 76), (15, 61, 78), (30, 56, 74), (43, 49, 68), (58, 51, 56), (53, 46, 70), (35, 41, 77), (32, 35, 78), (92, 59, 30), (136, 77, 0), (137, 73, 0), (141, 73, 0), (147, 76, 0), (155, 83, 12), (165, 92, 24), (170, 97, 31), (173, 101, 32), (176, 96, 20), (178, 91, 2), (178, 94, 0), (188, 99, 0), (193, 102, 0), (191, 100, 0), (187, 92, 3), (185, 86, 5), (181, 84, 1), (181, 83, 3), (198, 83, 19), (207, 75, 8), (221, 79, 2), (223, 80, 1), (223, 82, 1), (225, 84, 0), (227, 86, 0), (229, 89, 1), (230, 89, 0), (230, 89, 1), (230, 89, 0), (231, 90, 1), (231, 91, 1), (231, 91, 0), (232, 91, 1), (232, 91, 1), (232, 92, 1), (232, 91, 0), (232, 90, 0), (231, 91, 1), (229, 89, 0), (229, 87, 1), (230, 86, 1), (228, 83, 1), (226, 81, 0), (225, 79, 0), (223, 77, 0), (224, 76, 0), (223, 75, 1), (222, 73, 1), (221, 71, 0), (218, 69, 0), (217, 66, 1), (216, 64, 2), (214, 62, 2), (212, 60, 2), (211, 57, 2), (209, 55, 1), (208, 52, 2), (209, 48, 2), (208, 39, 0), (198, 36, 0), (178, 29, 3), (162, 4, 2), (153, 0, 3), (153, 2, 2), (152, 0, 1), (151, 1, 1), (151, 1, 1), (153, 1, 0), (154, 1, 0), (154, 1, 1), (154, 1, 1), (153, 1, 1), (151, 0, 2), (147, 1, 1), (145, 1, 1), (144, 1, 0), (142, 0, 0), (141, 0, 1), (138, 1, 1), (136, 0, 0), (137, 0, 1), (136, 1, 1), (135, 2, 2), (143, 1, 1), (150, 2, 1), (154, 3, 2), (159, 1, 2), (166, 3, 2), (173, 2, 3), (177, 1, 4), (165, 3, 7), (162, 2, 5), (165, 1, 3), (174, 1, 1), (185, 2, 3), (172, 216, 245), (171, 215, 248), (166, 213, 246), (162, 214, 243), (159, 213, 241), (156, 213, 243), (154, 210, 245), (153, 209, 246), (151, 208, 248), (151, 208, 245), (151, 207, 246), (147, 203, 244), (142, 203, 241), (141, 199, 243), (135, 202, 248), (54, 172, 206), (0, 129, 152), (0, 107, 115), (2, 90, 100), (0, 79, 86), (3, 80, 96), (23, 95, 137), (43, 117, 167), (52, 129, 187), (52, 130, 200), (45, 128, 199), (33, 117, 186), (22, 104, 154), (6, 85, 109), (0, 70, 75), (1, 67, 70), (0, 64, 65), (29, 101, 133), (67, 147, 217), (56, 132, 204), (36, 126, 198), (13, 124, 196), (1, 121, 196), (0, 120, 198), (3, 117, 195), (14, 113, 193), (27, 113, 195), (39, 110, 195), (47, 109, 195), (49, 112, 198), (51, 113, 200), (57, 114, 202), (69, 117, 206), (80, 120, 208), (89, 124, 210), (97, 131, 214), (106, 139, 216), (115, 144, 218), (128, 155, 227), (116, 151, 207), (10, 67, 86), (0, 59, 73), (5, 59, 76), (16, 58, 76), (37, 59, 77), (55, 52, 59), (41, 37, 50), (32, 36, 67), (37, 33, 68), (89, 50, 7), (118, 65, 0), (138, 86, 39), (171, 120, 106), (191, 145, 163), (197, 157, 202), (202, 167, 216), (195, 164, 214), (191, 161, 213), (200, 155, 207), (194, 139, 175), (189, 132, 130), (191, 114, 62), (186, 101, 11), (187, 98, 0), (190, 101, 0), (189, 98, 0), (185, 93, 0), (192, 98, 15), (185, 94, 17), (171, 69, 3), (189, 67, 10), (214, 78, 11), (222, 80, 1), (224, 82, 0), (225, 84, 2), (224, 84, 1), (224, 85, 0), (226, 86, 1), (226, 86, 0), (228, 87, 1), (228, 87, 1), (228, 87, 1), (229, 88, 2), (229, 88, 2), (228, 87, 2), (227, 86, 2), (226, 85, 0), (227, 86, 1), (226, 85, 1), (224, 82, 1), (225, 81, 1), (223, 79, 0), (222, 77, 0), (220, 75, 0), (218, 73, 0), (219, 72, 0), (219, 70, 0), (217, 68, 1), (214, 67, 1), (213, 64, 1), (212, 61, 1), (209, 59, 1), (207, 56, 2), (205, 54, 2), (204, 51, 1), (203, 47, 4), (202, 43, 1), (194, 32, 0), (196, 46, 37), (183, 77, 102), (137, 11, 15), (153, 0, 0), (152, 2, 2), (150, 1, 1), (149, 0, 1), (148, 0, 0), (148, 1, 1), (150, 1, 1), (151, 1, 1), (151, 1, 1), (151, 1, 1), (150, 1, 1), (147, 1, 3), (144, 2, 2), (143, 1, 2), (142, 0, 1), (140, 0, 0), (136, 2, 0), (131, 3, 0), (136, 0, 0), (140, 1, 1), (148, 1, 1), (152, 1, 0), (150, 0, 1), (145, 1, 0), (143, 1, 0), (143, 1, 0), (144, 1, 0), (147, 2, 0), (152, 2, 3), (110, 1, 2), (96, 4, 0), (143, 3, 1), (173, 0, 2), (182, 1, 3), (148, 206, 241), (143, 205, 240), (138, 202, 240), (136, 202, 241), (133, 200, 242), (130, 200, 243), (128, 198, 241), (126, 198, 240), (122, 198, 241), (124, 198, 240), (124, 196, 239), (118, 193, 238), (109, 189, 236), (96, 183, 236), (88, 175, 232), (83, 177, 233), (21, 149, 185), (0, 103, 113), (3, 89, 108), (30, 112, 158), (57, 140, 217), (63, 151, 248), (58, 149, 249), (51, 142, 246), (45, 139, 248), (40, 139, 251), (35, 142, 249), (29, 143, 249), (15, 133, 236), (11, 112, 181), (5, 78, 111), (1, 56, 55), (13, 83, 112), (28, 128, 212), (18, 121, 198), (8, 116, 189), (3, 114, 189), (1, 114, 190), (0, 111, 189), (1, 107, 186), (4, 103, 184), (9, 103, 184), (14, 104, 185), (25, 101, 185), (34, 100, 186), (41, 100, 190), (47, 101, 193), (61, 101, 197), (69, 104, 201), (76, 109, 204), (83, 115, 207), (92, 122, 209), (102, 132, 214), (111, 144, 224), (98, 133, 197), (4, 51, 73), (0, 49, 65), (4, 59, 78), (20, 65, 83), (30, 54, 75), (41, 40, 47), (56, 37, 30), (55, 32, 26), (52, 24, 20), (113, 72, 73), (178, 137, 164), (205, 174, 233), (214, 190, 255), (213, 188, 255), (206, 181, 248), (196, 171, 242), (187, 161, 233), (190, 162, 234), (190, 159, 234), (181, 149, 229), (183, 148, 233), (198, 157, 233), (197, 149, 183), (191, 122, 101), (186, 101, 16), (190, 102, 0), (189, 103, 3), (194, 106, 22), (175, 87, 3), (163, 72, 5), (109, 42, 10), (122, 42, 12), (200, 68, 8), (221, 76, 4), (221, 81, 2), (219, 80, 0), (219, 81, 0), (220, 82, 0), (222, 83, 0), (225, 83, 1), (225, 83, 3), (225, 83, 3), (225, 83, 1), (225, 83, 1), (225, 83, 2), (224, 82, 1), (223, 81, 0), (223, 82, 0), (222, 80, 0), (221, 78, 1), (221, 76, 1), (219, 75, 0), (218, 73, 0), (216, 71, 0), (212, 69, 1), (212, 68, 2), (211, 64, 1), (209, 61, 0), (207, 59, 1), (204, 57, 1), (203, 53, 1), (202, 51, 0), (202, 50, 0), (201, 48, 0), (202, 44, 0), (198, 37, 0), (182, 37, 16), (180, 65, 106), (195, 129, 222), (186, 103, 168), (147, 1, 8), (150, 1, 0), (148, 1, 2), (147, 1, 2), (146, 0, 2), (145, 0, 1), (146, 1, 0), (146, 1, 0), (148, 2, 1), (147, 1, 1), (147, 1, 1), (146, 2, 1), (144, 2, 2), (142, 1, 1), (141, 1, 0), (139, 1, 0), (137, 0, 0), (132, 2, 0), (133, 2, 0), (149, 0, 1), (156, 0, 2), (158, 0, 0), (161, 0, 0), (160, 1, 0), (156, 1, 0), (156, 0, 1), (156, 0, 1), (154, 1, 1), (152, 1, 1), (148, 1, 1), (138, 3, 2), (119, 3, 1), (149, 3, 2), (175, 1, 2), (178, 2, 2), (123, 192, 234), (115, 188, 231), (108, 187, 233), (104, 186, 237), (103, 185, 236), (99, 187, 236), (96, 186, 234), (95, 185, 234), (94, 185, 234), (94, 185, 234), (91, 182, 234), (74, 178, 230), (65, 175, 232), (48, 164, 224), (45, 160, 221), (42, 152, 215), (18, 148, 197), (13, 117, 151), (43, 137, 198), (41, 148, 240), (22, 134, 241), (8, 124, 235), (3, 120, 233), (2, 118, 232), (2, 118, 231), (3, 119, 233), (2, 120, 233), (0, 123, 233), (0, 130, 238), (5, 136, 243), (11, 130, 222), (10, 86, 131), (3, 66, 90), (5, 111, 195), (0, 112, 193), (1, 109, 186), (2, 110, 185), (3, 109, 185), (0, 104, 181), (0, 101, 179), (1, 100, 180), (0, 98, 178), (0, 96, 177), (5, 92, 177), (15, 92, 180), (22, 91, 183), (30, 91, 185), (45, 91, 191), (53, 93, 194), (60, 100, 198), (68, 103, 198), (77, 107, 199), (88, 119, 207), (95, 130, 216), (69, 140, 202), (8, 118, 138), (7, 70, 98), (9, 55, 78), (9, 54, 71), (24, 41, 65), (40, 34, 42), (51, 23, 15), (68, 38, 37), (143, 114, 156), (199, 172, 243), (207, 176, 255), (197, 167, 247), (190, 161, 237), (188, 159, 233), (184, 151, 228), (179, 143, 227), (176, 138, 226), (177, 136, 225), (176, 134, 222), (175, 131, 216), (173, 128, 211), (178, 133, 217), (189, 146, 232), (200, 153, 245), (197, 142, 185), (184, 109, 58), (185, 101, 12), (185, 102, 11), (168, 80, 0), (161, 69, 5), (80, 33, 8), (73, 7, 4), (138, 11, 4), (158, 25, 6), (188, 58, 6), (213, 75, 8), (218, 76, 5), (216, 77, 0), (217, 79, 0), (220, 79, 0), (222, 79, 3), (220, 78, 4), (219, 78, 2), (221, 78, 2), (220, 77, 1), (219, 77, 0), (220, 77, 1), (219, 76, 1), (218, 75, 1), (217, 74, 1), (217, 74, 2), (215, 71, 1), (214, 70, 1), (212, 68, 1), (210, 65, 1), (208, 63, 2), (205, 59, 1), (203, 56, 1), (203, 54, 2), (201, 51, 2), (201, 50, 1), (200, 49, 1), (198, 47, 0), (192, 44, 0), (173, 38, 23), (163, 46, 82), (165, 75, 164), (165, 101, 217), (166, 106, 215), (148, 26, 48), (146, 0, 0), (147, 1, 3), (145, 0, 2), (144, 0, 1), (144, 0, 1), (144, 0, 1), (146, 0, 1), (146, 0, 2), (146, 1, 2), (146, 0, 2), (146, 0, 2), (146, 0, 1), (144, 0, 1), (142, 0, 0), (141, 0, 0), (139, 0, 1), (135, 1, 0), (131, 2, 1), (141, 2, 1), (161, 0, 3), (164, 0, 3), (162, 1, 0), (163, 1, 0), (163, 1, 0), (164, 0, 0), (164, 0, 1), (164, 0, 2), (162, 0, 1), (158, 0, 1), (153, 2, 1), (148, 2, 1), (146, 1, 1), (155, 2, 1), (174, 3, 0), (175, 1, 1), (88, 174, 229), (75, 172, 228), (63, 172, 229), (59, 170, 229), (61, 171, 230), (55, 173, 232), (51, 172, 232), (51, 172, 232), (53, 171, 232), (51, 171, 231), (40, 168, 228), (26, 164, 228), (19, 158, 227), (3, 148, 217), (1, 148, 215), (0, 130, 200), (10, 131, 201), (35, 149, 231), (20, 131, 241), (0, 115, 231), (1, 112, 228), (0, 109, 225), (0, 107, 225), (0, 106, 227), (0, 107, 228), (0, 107, 229), (0, 108, 229), (0, 108, 229), (2, 112, 228), (4, 118, 225), (1, 124, 229), (6, 125, 223), (7, 82, 139), (8, 84, 161), (2, 104, 195), (1, 104, 184), (2, 105, 183), (1, 104, 181), (0, 100, 177), (0, 97, 174), (1, 97, 175), (0, 95, 175), (1, 93, 177), (1, 91, 180), (1, 88, 180), (3, 87, 178), (8, 86, 178), (19, 88, 185), (21, 88, 186), (24, 91, 188), (42, 95, 192), (59, 104, 200), (72, 111, 206), (71, 122, 207), (30, 157, 209), (6, 190, 214), (10, 170, 203), (6, 87, 115), (10, 34, 52), (31, 34, 45), (28, 18, 20), (68, 45, 70), (172, 141, 208), (204, 171, 255), (190, 157, 246), (182, 149, 235), (178, 140, 232), (171, 132, 227), (165, 125, 223), (161, 117, 219), (157, 110, 214), (154, 106, 207), (155, 105, 207), (147, 96, 201), (151, 94, 199), (165, 107, 208), (163, 108, 203), (167, 114, 205), (176, 126, 217), (187, 139, 236), (197, 144, 220), (190, 122, 117), (163, 81, 7), (157, 72, 0), (145, 55, 4), (71, 19, 6), (81, 4, 9), (112, 6, 11), (106, 3, 11), (125, 20, 20), (138, 30, 11), (163, 52, 22), (188, 65, 19), (202, 68, 5), (215, 78, 6), (222, 78, 2), (217, 76, 1), (216, 75, 2), (214, 74, 1), (213, 75, 0), (214, 75, 0), (214, 75, 1), (213, 73, 0), (212, 72, 1), (212, 70, 3), (212, 69, 2), (210, 67, 1), (208, 65, 1), (207, 64, 1), (206, 61, 0), (202, 56, 0), (199, 52, 0), (197, 49, 0), (199, 48, 0), (195, 45, 0), (188, 46, 0), (176, 42, 11), (160, 37, 44), (139, 40, 90), (130, 47, 147), (131, 60, 177), (135, 63, 176), (142, 67, 185), (145, 53, 133), (143, 2, 6), (147, 2, 0), (145, 0, 2), (144, 0, 0), (142, 0, 0), (142, 0, 0), (142, 0, 0), (143, 0, 0), (144, 1, 1), (144, 1, 0), (144, 1, 1), (144, 1, 1), (144, 1, 0), (143, 0, 0), (140, 0, 0), (138, 0, 0), (135, 0, 2), (132, 1, 1), (135, 0, 1), (150, 2, 2), (160, 1, 2), (161, 0, 2), (161, 1, 1), (163, 0, 0), (164, 0, 0), (163, 0, 0), (163, 1, 0), (162, 1, 0), (161, 1, 0), (158, 0, 1), (154, 1, 1), (149, 1, 1), (144, 0, 1), (152, 2, 0), (165, 0, 0), (167, 0, 0), (43, 157, 212), (16, 153, 212), (4, 153, 216), (7, 155, 216), (13, 157, 220), (7, 155, 220), (0, 154, 219), (0, 151, 220), (0, 154, 224), (2, 156, 226), (2, 154, 221), (2, 150, 222), (2, 146, 219), (1, 139, 214), (0, 130, 205), (7, 123, 200), (23, 140, 221), (9, 126, 226), (0, 110, 227), (0, 102, 223), (1, 97, 217), (0, 93, 215), (0, 93, 217), (0, 93, 222), (1, 92, 222), (1, 92, 223), (2, 93, 224), (2, 94, 223), (1, 98, 220), (1, 104, 219), (3, 107, 220), (1, 109, 220), (6, 94, 198), (5, 62, 155), (2, 90, 176), (0, 99, 181), (2, 101, 180), (1, 102, 177), (0, 99, 174), (0, 97, 173), (0, 97, 174), (1, 95, 175), (1, 93, 176), (0, 91, 179), (0, 89, 179), (0, 87, 178), (1, 85, 179), (2, 84, 181), (0, 84, 183), (1, 85, 184), (13, 88, 188), (28, 97, 196), (43, 106, 204), (38, 122, 202), (9, 156, 199), (0, 174, 204), (0, 179, 207), (8, 166, 198), (15, 62, 88), (20, 12, 17), (63, 47, 82), (174, 146, 226), (191, 159, 253), (178, 143, 236), (171, 131, 228), (163, 122, 219), (155, 114, 214), (148, 105, 209), (143, 96, 203), (137, 86, 197), (132, 80, 190), (128, 76, 182), (127, 74, 178), (127, 72, 175), (131, 74, 178), (139, 79, 183), (140, 80, 180), (145, 83, 183), (155, 90, 189), (164, 101, 196), (177, 125, 215), (198, 149, 227), (178, 108, 130), (132, 59, 20), (122, 49, 33), (97, 39, 56), (99, 33, 57), (98, 23, 47), (90, 8, 33), (89, 3, 31), (80, 4, 18), (81, 11, 16), (89, 14, 13), (104, 18, 7), (137, 31, 10), (167, 48, 6), (192, 60, 4), (206, 65, 6), (212, 69, 3), (208, 70, 0), (209, 69, 0), (211, 70, 0), (210, 69, 0), (208, 67, 0), (209, 64, 3), (208, 62, 2), (206, 60, 0), (203, 60, 0), (202, 58, 0), (203, 55, 1), (203, 52, 2), (197, 49, 3), (189, 46, 1), (176, 42, 5), (166, 47, 35), (131, 30, 62), (109, 22, 90), (101, 26, 123), (100, 29, 132), (104, 31, 131), (106, 30, 130), (103, 30, 132), (108, 38, 141), (124, 14, 60), (143, 0, 0), (144, 0, 0), (146, 0, 1), (145, 0, 1), (142, 0, 0), (141, 0, 0), (141, 0, 0), (141, 0, 0), (141, 0, 0), (141, 1, 0), (141, 1, 0), (141, 1, 0), (141, 1, 0), (140, 0, 0), (138, 0, 1), (136, 0, 1), (134, 0, 1), (130, 1, 0), (136, 1, 1), (149, 1, 2), (152, 1, 1), (152, 1, 1), (152, 2, 1), (154, 2, 0), (158, 2, 1), (160, 1, 1), (161, 1, 1), (160, 1, 1), (159, 1, 0), (156, 1, 1), (153, 1, 0), (149, 1, 1), (140, 0, 0), (151, 1, 0), (194, 33, 30), (228, 77, 73), (49, 157, 207), (92, 188, 222), (132, 208, 235), (159, 220, 240), (167, 225, 244), (164, 222, 243), (139, 215, 234), (95, 193, 227), (49, 164, 221), (4, 141, 209), (0, 138, 213), (1, 141, 213), (2, 136, 209), (1, 129, 206), (1, 119, 197), (15, 131, 214), (9, 123, 225), (0, 105, 217), (0, 96, 216), (1, 88, 213), (0, 86, 209), (0, 84, 207), (0, 82, 208), (0, 83, 209), (1, 85, 208), (0, 86, 208), (1, 87, 209), (2, 88, 211), (2, 89, 212), (0, 92, 212), (1, 96, 213), (1, 95, 208), (1, 84, 195), (0, 52, 148), (4, 56, 145), (3, 90, 177), (0, 98, 177), (1, 100, 175), (0, 99, 171), (1, 99, 172), (2, 99, 175), (2, 97, 178), (2, 95, 178), (1, 94, 180), (0, 91, 180), (0, 89, 180), (2, 85, 181), (1, 83, 182), (0, 84, 185), (1, 86, 189), (0, 91, 190), (2, 98, 195), (8, 107, 197), (5, 119, 188), (0, 145, 187), (0, 159, 193), (0, 162, 196), (1, 166, 201), (8, 110, 139), (40, 46, 79), (160, 137, 216), (184, 152, 248), (170, 132, 227), (160, 120, 220), (150, 107, 211), (141, 97, 204), (135, 89, 198), (128, 80, 190), (120, 72, 182), (114, 63, 175), (109, 57, 168), (105, 53, 162), (104, 50, 155), (102, 48, 148), (105, 50, 147), (109, 52, 147), (117, 56, 151), (125, 61, 158), (130, 62, 162), (136, 67, 164), (156, 91, 183), (163, 102, 187), (155, 92, 164), (122, 59, 102), (114, 54, 97), (99, 42, 84), (89, 33, 72), (83, 25, 62), (82, 14, 50), (81, 1, 40), (79, 0, 34), (77, 0, 28), (79, 2, 18), (79, 2, 16), (78, 0, 16), (81, 4, 9), (98, 12, 5), (117, 15, 6), (144, 24, 10), (169, 37, 23), (177, 37, 24), (183, 40, 9), (185, 45, 6), (186, 47, 5), (189, 47, 3), (187, 48, 1), (183, 43, 9), (175, 39, 12), (169, 37, 12), (158, 33, 12), (146, 24, 12), (126, 9, 16), (109, 0, 21), (109, 8, 48), (138, 60, 113), (138, 75, 148), (138, 79, 152), (150, 99, 163), (163, 111, 174), (171, 120, 185), (172, 120, 186), (165, 112, 179), (153, 102, 167), (158, 71, 108), (160, 33, 44), (141, 6, 12), (132, 0, 0), (137, 0, 0), (143, 0, 0), (142, 0, 0), (141, 0, 0), (141, 0, 0), (141, 0, 0), (141, 0, 0), (141, 0, 0), (141, 0, 0), (139, 0, 0), (139, 0, 1), (138, 1, 2), (137, 1, 1), (134, 1, 0), (130, 1, 0), (133, 1, 2), (141, 1, 2), (143, 0, 0), (144, 0, 1), (146, 1, 1), (147, 1, 1), (150, 1, 1), (154, 0, 1), (154, 1, 0), (154, 1, 0), (153, 1, 0), (153, 1, 0), (150, 1, 1), (141, 0, 0), (156, 13, 15), (220, 70, 65), (255, 100, 85), (255, 100, 82), (196, 235, 245), (217, 246, 255), (215, 242, 255), (215, 241, 254), (220, 242, 254), (218, 243, 255), (219, 246, 255), (219, 245, 254), (207, 237, 249), (147, 214, 239), (53, 165, 211), (0, 123, 203), (0, 125, 207), (2, 122, 202), (3, 121, 205), (6, 119, 220), (2, 97, 208), (1, 85, 200), (0, 82, 199), (1, 79, 198), (0, 76, 198), (2, 74, 199), (3, 73, 199), (3, 74, 197), (1, 75, 196), (1, 75, 199), (1, 75, 198), (1, 76, 199), (1, 77, 202), (0, 81, 201), (2, 83, 198), (1, 81, 193), (1, 75, 183), (2, 56, 154), (2, 32, 112), (4, 63, 146), (1, 89, 175), (1, 96, 173), (1, 97, 170), (1, 100, 173), (2, 101, 177), (2, 100, 180), (2, 98, 182), (2, 96, 182), (2, 93, 183), (1, 91, 183), (2, 87, 184), (1, 85, 184), (1, 86, 186), (1, 89, 191), (0, 94, 196), (0, 103, 205), (0, 102, 174), (0, 97, 146), (0, 117, 160), (0, 135, 175), (0, 141, 186), (1, 143, 180), (61, 183, 200), (157, 165, 224), (176, 136, 240), (162, 122, 228), (151, 109, 214), (141, 96, 205), (132, 85, 197), (124, 77, 191), (118, 68, 182), (107, 57, 169), (98, 50, 159), (93, 46, 149), (93, 43, 142), (92, 40, 136), (90, 38, 131), (88, 35, 127), (87, 35, 121), (86, 33, 116), (92, 35, 119), (100, 40, 124), (96, 35, 121), (111, 51, 132), (148, 87, 163), (145, 79, 155), (128, 63, 134), (114, 54, 122), (102, 46, 105), (91, 37, 88), (84, 30, 75), (78, 26, 63), (73, 20, 54), (70, 9, 45), (71, 2, 38), (72, 0, 34), (75, 0, 31), (77, 1, 24), (78, 2, 23), (79, 1, 25), (80, 1, 16), (79, 2, 5), (84, 1, 13), (124, 11, 57), (133, 2, 67), (126, 0, 51), (124, 1, 37), (124, 2, 33), (127, 3, 29), (132, 4, 32), (120, 5, 37), (95, 4, 30), (88, 0, 20), (77, 0, 5), (73, 0, 8), (95, 17, 59), (139, 69, 118), (182, 125, 169), (205, 163, 205), (212, 184, 224), (219, 195, 235), (222, 199, 237), (225, 201, 239), (225, 201, 239), (227, 203, 240), (230, 204, 242), (231, 203, 242), (229, 202, 239), (221, 196, 232), (211, 172, 202), (195, 127, 152), (165, 68, 86), (140, 10, 16), (131, 0, 0), (138, 0, 0), (141, 0, 0), (141, 0, 0), (141, 0, 0), (141, 0, 0), (141, 0, 0), (139, 0, 1), (139, 0, 3), (138, 1, 2), (136, 1, 1), (133, 1, 1), (130, 1, 1), (128, 0, 2), (130, 1, 1), (133, 1, 0), (135, 0, 0), (137, 1, 1), (139, 1, 0), (143, 1, 0), (144, 1, 0), (145, 1, 0), (144, 2, 0), (145, 1, 0), (148, 0, 1), (141, 0, 0), (160, 15, 15), (237, 76, 64), (252, 88, 68), (243, 82, 63), (247, 76, 57), (195, 228, 247), (194, 231, 254), (192, 230, 251), (187, 229, 248), (189, 230, 247), (191, 231, 250), (192, 230, 252), (192, 231, 253), (191, 232, 253), (200, 237, 254), (191, 236, 255), (106, 184, 231), (9, 119, 198), (0, 113, 199), (4, 119, 209), (1, 100, 204), (4, 82, 197), (2, 76, 191), (1, 73, 188), (1, 70, 187), (0, 68, 189), (1, 67, 189), (3, 65, 189), (3, 64, 188), (2, 64, 189), (1, 65, 191), (1, 67, 192), (2, 68, 193), (1, 68, 193), (0, 70, 190), (2, 71, 185), (3, 72, 182), (2, 69, 178), (3, 57, 159), (2, 33, 111), (0, 38, 88), (2, 67, 139), (3, 81, 165), (4, 89, 165), (2, 94, 170), (0, 98, 178), (1, 99, 181), (1, 98, 182), (1, 95, 182), (1, 93, 184), (1, 91, 184), (2, 89, 185), (0, 88, 186), (0, 88, 189), (0, 90, 196), (0, 86, 193), (6, 91, 180), (46, 107, 157), (82, 135, 167), (80, 150, 178), (53, 146, 172), (8, 124, 162), (28, 175, 194), (135, 197, 240), (170, 130, 226), (160, 114, 222), (142, 99, 211), (132, 87, 199), (127, 79, 192), (121, 70, 186), (109, 59, 173), (99, 49, 161), (92, 43, 150), (87, 39, 143), (84, 36, 132), (81, 32, 124), (80, 29, 116), (77, 28, 111), (75, 25, 108), (72, 21, 102), (74, 21, 99), (77, 21, 99), (75, 19, 92), (83, 27, 100), (151, 95, 169), (166, 108, 184), (145, 83, 162), (127, 66, 140), (107, 50, 116), (93, 38, 99), (84, 31, 88), (78, 25, 76), (71, 22, 63), (65, 19, 53), (60, 13, 47), (59, 7, 41), (61, 2, 37), (63, 0, 32), (65, 1, 27), (67, 0, 25), (71, 1, 24), (76, 0, 19), (79, 1, 14), (79, 1, 13), (85, 0, 17), (106, 2, 33), (117, 4, 56), (113, 2, 58), (112, 2, 51), (115, 2, 52), (109, 2, 45), (83, 2, 25), (67, 0, 12), (58, 0, 0), (94, 30, 43), (158, 102, 124), (199, 160, 202), (220, 187, 234), (221, 195, 241), (217, 196, 235), (214, 197, 234), (213, 197, 234), (213, 195, 233), (214, 196, 233), (217, 199, 235), (219, 200, 237), (219, 201, 238), (218, 202, 238), (220, 201, 239), (219, 205, 242), (224, 214, 247), (234, 218, 253), (233, 211, 247), (222, 173, 207), (181, 102, 116), (141, 19, 21), (131, 0, 0), (141, 0, 0), (142, 0, 1), (139, 0, 1), (139, 0, 2), (139, 0, 2), (138, 1, 4), (137, 0, 2), (134, 0, 2), (132, 1, 2), (130, 1, 1), (127, 1, 0), (126, 1, 0), (128, 1, 0), (130, 1, 1), (133, 1, 2), (136, 0, 1), (138, 0, 0), (139, 0, 0), (139, 0, 0), (138, 1, 0), (139, 0, 0), (138, 0, 1), (140, 4, 4), (222, 61, 56), (246, 72, 54), (237, 63, 42), (236, 61, 43), (235, 58, 41), (177, 222, 250), (175, 222, 250), (171, 221, 248), (167, 221, 246), (170, 222, 249), (173, 223, 250), (174, 223, 250), (172, 223, 251), (170, 223, 251), (170, 222, 251), (173, 221, 250), (181, 227, 253), (110, 189, 236), (10, 112, 193), (2, 106, 199), (1, 86, 191), (4, 72, 186), (1, 68, 183), (0, 65, 181), (0, 62, 181), (0, 61, 181), (0, 60, 180), (1, 59, 180), (1, 59, 180), (1, 59, 180), (1, 59, 181), (0, 60, 181), (0, 61, 181), (0, 62, 182), (0, 61, 178), (0, 64, 176), (1, 64, 174), (0, 63, 168), (1, 53, 153), (1, 35, 121), (0, 38, 64), (1, 51, 77), (3, 56, 119), (3, 57, 132), (3, 63, 140), (0, 70, 148), (1, 76, 159), (2, 83, 169), (3, 88, 176), (2, 87, 178), (0, 88, 182), (1, 88, 184), (1, 88, 186), (0, 83, 190), (0, 79, 179), (91, 142, 198), (191, 201, 227), (233, 225, 243), (247, 232, 251), (245, 230, 251), (234, 227, 246), (201, 211, 228), (150, 213, 226), (140, 137, 215), (149, 98, 217), (136, 91, 206), (124, 77, 192), (118, 71, 186), (112, 65, 179), (102, 54, 166), (93, 44, 152), (87, 38, 141), (79, 32, 132), (75, 30, 125), (74, 27, 118), (73, 22, 111), (69, 18, 105), (66, 17, 98), (64, 15, 93), (63, 11, 88), (64, 9, 85), (60, 6, 79), (67, 16, 88), (152, 101, 179), (172, 120, 205), (146, 93, 178), (128, 72, 157), (113, 60, 137), (96, 45, 114), (84, 34, 97), (76, 28, 85), (70, 23, 76), (65, 21, 65), (62, 19, 57), (60, 15, 52), (57, 11, 46), (55, 8, 42), (54, 5, 39), (54, 3, 37), (56, 1, 35), (58, 1, 32), (63, 2, 29), (67, 1, 25), (71, 2, 21), (75, 2, 20), (81, 0, 16), (96, 2, 30), (114, 2, 57), (116, 1, 65), (107, 3, 56), (74, 1, 31), (46, 0, 7), (70, 13, 25), (143, 95, 123), (204, 167, 214), (215, 188, 233), (208, 188, 233), (209, 186, 229), (212, 188, 231), (211, 190, 231), (211, 192, 233), (212, 191, 234), (211, 190, 234), (212, 193, 234), (214, 195, 234), (214, 196, 235), (215, 197, 236), (215, 197, 238), (215, 198, 238), (218, 201, 238), (221, 203, 237), (223, 205, 238), (221, 205, 237), (223, 214, 244), (233, 222, 253), (224, 185, 219), (173, 88, 101), (136, 1, 1), (136, 0, 0), (137, 2, 3), (138, 1, 3), (139, 0, 2), (138, 1, 2), (137, 0, 0), (135, 0, 0), (133, 1, 1), (130, 1, 1), (127, 1, 0), (126, 1, 0), (126, 1, 1), (126, 1, 2), (129, 2, 2), (130, 1, 0), (132, 0, 0), (134, 0, 0), (135, 0, 2), (135, 0, 1), (135, 1, 1), (125, 0, 0), (173, 32, 30), (234, 67, 54), (231, 52, 27), (230, 48, 24), (229, 44, 18), (228, 43, 14), (152, 213, 244), (154, 212, 243), (154, 212, 243), (154, 213, 245), (155, 214, 245), (156, 215, 245), (156, 215, 245), (156, 215, 245), (156, 213, 246), (155, 213, 248), (147, 210, 246), (141, 206, 243), (146, 212, 243), (81, 169, 226), (3, 90, 192), (2, 71, 181), (4, 65, 176), (2, 61, 173), (0, 57, 173), (0, 55, 173), (1, 55, 173), (0, 54, 172), (1, 54, 171), (1, 54, 171), (1, 54, 172), (2, 54, 173), (1, 54, 172), (1, 55, 172), (0, 56, 172), (0, 57, 170), (0, 58, 169), (0, 58, 169), (1, 58, 160), (1, 51, 145), (1, 34, 127), (5, 44, 93), (2, 59, 83), (2, 57, 88), (3, 57, 102), (3, 57, 104), (1, 50, 100), (1, 45, 105), (2, 48, 124), (5, 60, 152), (7, 68, 164), (2, 71, 169), (1, 72, 171), (0, 67, 171), (11, 66, 161), (144, 169, 208), (245, 232, 254), (237, 215, 246), (226, 203, 247), (222, 202, 246), (224, 200, 242), (226, 202, 242), (237, 210, 246), (242, 217, 247), (223, 196, 237), (143, 107, 197), (110, 64, 184), (112, 64, 178), (106, 57, 172), (95, 49, 160), (87, 41, 148), (82, 35, 137), (76, 29, 126), (70, 24, 118), (67, 21, 113), (64, 18, 103), (62, 14, 98), (59, 10, 93), (57, 8, 86), (58, 5, 81), (57, 4, 77), (55, 1, 72), (50, 0, 74), (134, 86, 170), (169, 121, 211), (142, 93, 183), (123, 75, 159), (109, 61, 142), (97, 49, 124), (85, 38, 107), (79, 32, 97), (72, 27, 86), (68, 23, 78), (65, 22, 70), (63, 19, 63), (60, 16, 56), (56, 14, 50), (55, 13, 46), (56, 10, 44), (55, 8, 42), (55, 6, 39), (56, 4, 35), (60, 2, 34), (65, 2, 32), (66, 0, 29), (70, 0, 28), (76, 1, 23), (81, 1, 15), (94, 1, 36), (107, 3, 68), (80, 1, 48), (42, 0, 17), (88, 43, 73), (184, 140, 178), (213, 181, 226), (206, 180, 224), (205, 179, 223), (205, 182, 225), (205, 184, 227), (207, 185, 228), (206, 187, 229), (206, 186, 231), (206, 185, 232), (208, 186, 234), (208, 184, 235), (207, 183, 234), (206, 187, 234), (208, 188, 237), (209, 188, 235), (209, 190, 235), (212, 193, 236), (215, 196, 236), (218, 200, 237), (217, 203, 236), (220, 205, 236), (223, 207, 238), (228, 214, 250), (235, 218, 250), (205, 151, 168), (141, 26, 33), (132, 0, 0), (141, 0, 1), (140, 0, 2), (138, 1, 3), (137, 1, 2), (137, 0, 1), (135, 0, 1), (133, 0, 2), (130, 0, 1), (128, 0, 0), (126, 1, 1), (125, 1, 3), (126, 1, 2), (128, 1, 1), (131, 1, 1), (132, 0, 1), (134, 0, 2), (134, 0, 2), (133, 1, 1), (135, 3, 4), (209, 44, 33), (226, 45, 17), (223, 35, 2), (221, 29, 1), (220, 26, 0), (221, 21, 0), (124, 199, 245), (125, 200, 245), (126, 201, 245), (127, 202, 247), (129, 204, 247), (131, 205, 248), (131, 205, 248), (132, 204, 246), (133, 202, 244), (129, 202, 244), (122, 199, 242), (113, 194, 238), (102, 188, 231), (81, 173, 230), (4, 86, 183), (0, 63, 169), (1, 60, 167), (0, 57, 164), (0, 54, 164), (0, 52, 163), (0, 50, 162), (0, 50, 161), (1, 50, 162), (1, 51, 163), (1, 50, 163), (1, 51, 163), (0, 51, 163), (0, 51, 163), (1, 52, 162), (0, 54, 162), (0, 55, 162), (0, 56, 162), (1, 56, 154), (3, 52, 141), (0, 34, 118), (4, 47, 105), (8, 114, 149), (5, 139, 168), (6, 139, 172), (3, 133, 167), (3, 117, 151), (1, 91, 129), (4, 61, 112), (1, 41, 113), (2, 42, 122), (2, 48, 131), (0, 53, 138), (2, 52, 134), (139, 159, 209), (237, 219, 248), (214, 185, 232), (204, 176, 231), (202, 174, 233), (203, 172, 233), (205, 173, 234), (207, 175, 235), (209, 178, 235), (213, 181, 235), (227, 198, 242), (215, 184, 234), (118, 73, 178), (95, 45, 161), (94, 45, 155), (84, 37, 143), (79, 33, 132), (72, 27, 122), (65, 21, 113), (62, 18, 108), (60, 15, 103), (56, 11, 94), (55, 8, 90), (52, 3, 83), (53, 2, 77), (53, 2, 74), (52, 1, 70), (42, 0, 58), (103, 53, 133), (169, 123, 215), (140, 93, 187), (122, 75, 168), (105, 61, 146), (98, 54, 134), (84, 41, 115), (78, 34, 104), (72, 28, 96), (69, 27, 87), (67, 25, 81), (64, 23, 74), (62, 21, 68), (59, 19, 62), (56, 17, 55), (56, 15, 51), (56, 15, 48), (57, 13, 45), (56, 11, 42), (55, 7, 40), (57, 4, 39), (61, 4, 38), (61, 0, 32), (61, 0, 28), (67, 2, 25), (73, 2, 18), (74, 1, 21), (84, 2, 36), (50, 0, 28), (106, 67, 95), (197, 160, 200), (205, 176, 223), (201, 173, 220), (201, 176, 219), (202, 176, 220), (200, 178, 222), (200, 179, 225), (202, 181, 227), (202, 181, 228), (202, 180, 228), (202, 181, 229), (203, 182, 230), (204, 180, 231), (203, 180, 230), (204, 182, 230), (206, 183, 232), (206, 183, 232), (208, 184, 233), (209, 186, 234), (210, 190, 234), (211, 194, 235), (214, 198, 237), (218, 200, 237), (221, 204, 238), (223, 207, 234), (226, 209, 237), (236, 219, 252), (221, 182, 215), (155, 53, 70), (133, 0, 0), (140, 1, 2), (138, 1, 4), (138, 1, 4), (138, 0, 3), (137, 0, 2), (136, 0, 1), (135, 1, 1), (132, 1, 1), (127, 1, 0), (124, 0, 1), (124, 0, 1), (128, 0, 1), (131, 2, 2), (132, 1, 2), (131, 1, 1), (132, 1, 1), (128, 0, 2), (145, 9, 10), (218, 38, 20), (218, 17, 1), (216, 8, 1), (219, 4, 0), (216, 0, 0), (208, 11, 7), (96, 187, 239), (97, 189, 238), (98, 190, 237), (99, 192, 239), (101, 194, 240), (104, 194, 241), (106, 193, 241), (106, 192, 241), (104, 191, 239), (98, 190, 238), (92, 187, 236), (85, 180, 234), (65, 175, 229), (34, 152, 216), (0, 82, 175), (1, 61, 163), (2, 57, 160), (1, 53, 157), (2, 50, 156), (1, 48, 152), (1, 46, 151), (2, 45, 151), (2, 46, 152), (2, 46, 152), (2, 46, 151), (2, 48, 150), (1, 48, 151), (1, 48, 152), (2, 48, 155), (1, 51, 156), (0, 53, 155), (2, 54, 156), (2, 54, 150), (3, 48, 135), (3, 39, 111), (7, 119, 160), (6, 166, 197), (3, 163, 195), (2, 159, 193), (0, 160, 192), (2, 153, 186), (4, 141, 175), (7, 124, 160), (4, 89, 137), (1, 45, 110), (3, 40, 111), (0, 46, 124), (58, 108, 168), (218, 205, 241), (200, 167, 227), (189, 153, 222), (187, 149, 221), (188, 148, 219), (189, 146, 219), (190, 147, 222), (194, 151, 225), (197, 154, 224), (197, 155, 223), (201, 159, 226), (218, 177, 235), (180, 134, 209), (83, 33, 142), (81, 33, 138), (75, 30, 127), (65, 21, 112), (57, 13, 102), (51, 7, 94), (51, 6, 93), (52, 9, 92), (50, 7, 86), (49, 3, 81), (48, 0, 76), (49, 0, 71), (48, 0, 68), (42, 0, 61), (60, 15, 83), (156, 112, 197), (144, 101, 199), (121, 76, 173), (107, 62, 156), (93, 52, 139), (85, 43, 125), (78, 35, 112), (73, 32, 104), (69, 28, 96), (65, 26, 88), (64, 25, 82), (61, 23, 76), (59, 21, 72), (58, 21, 67), (55, 19, 60), (54, 18, 57), (54, 17, 53), (56, 15, 50), (56, 13, 47), (53, 11, 45), (56, 11, 46), (54, 5, 40), (54, 3, 34), (57, 2, 31), (62, 2, 29), (69, 2, 24), (74, 0, 19), (67, 0, 12), (118, 75, 105), (197, 165, 208), (198, 168, 214), (195, 166, 214), (195, 169, 216), (194, 171, 216), (194, 172, 218), (194, 173, 219), (196, 174, 222), (197, 175, 224), (196, 174, 225), (196, 174, 224), (196, 174, 223), (197, 175, 224), (198, 174, 226), (198, 174, 226), (199, 175, 227), (202, 176, 229), (202, 176, 228), (204, 179, 229), (206, 181, 232), (206, 183, 233), (207, 187, 232), (212, 193, 235), (216, 197, 237), (219, 201, 237), (221, 205, 235), (224, 207, 237), (225, 207, 239), (229, 212, 247), (230, 197, 228), (158, 69, 80), (126, 0, 0), (139, 0, 2), (139, 0, 4), (139, 0, 3), (137, 0, 0), (137, 0, 0), (138, 1, 0), (135, 1, 1), (132, 1, 1), (128, 0, 0), (126, 0, 0), (126, 1, 1), (127, 2, 1), (129, 1, 1), (129, 1, 1), (128, 2, 2), (122, 1, 2), (146, 10, 9), (214, 17, 8), (212, 0, 0), (208, 0, 0), (203, 0, 0), (220, 33, 29), (247, 89, 78), (56, 178, 229), (59, 178, 232), (62, 178, 235), (65, 180, 236), (69, 181, 235), (71, 181, 233), (71, 182, 234), (73, 180, 234), (72, 179, 235), (64, 176, 235), (54, 171, 232), (42, 163, 226), (16, 159, 218), (7, 143, 208), (1, 84, 173), (3, 60, 159), (2, 55, 155), (1, 52, 151), (2, 49, 148), (1, 47, 143), (1, 47, 142), (0, 46, 142), (1, 45, 144), (2, 44, 145), (2, 44, 144), (3, 45, 143), (4, 46, 145), (4, 46, 146), (2, 47, 146), (1, 50, 147), (0, 52, 150), (2, 52, 152), (2, 52, 144), (1, 41, 123), (10, 89, 143), (4, 167, 189), (2, 158, 185), (2, 156, 186), (0, 153, 186), (0, 151, 185), (1, 148, 183), (0, 146, 178), (1, 141, 174), (3, 132, 170), (6, 87, 143), (0, 40, 112), (0, 57, 131), (146, 159, 212), (199, 164, 222), (171, 131, 209), (169, 126, 204), (169, 123, 203), (170, 122, 203), (175, 123, 206), (178, 124, 210), (180, 127, 211), (182, 130, 210), (183, 131, 207), (185, 134, 211), (189, 135, 211), (199, 147, 217), (105, 56, 150), (59, 14, 117), (59, 17, 110), (78, 37, 124), (93, 51, 136), (93, 48, 133), (76, 29, 112), (46, 1, 80), (39, 0, 70), (47, 2, 77), (46, 0, 73), (44, 0, 68), (44, 0, 64), (35, 0, 56), (110, 67, 142), (158, 113, 207), (125, 79, 182), (108, 63, 161), (96, 51, 148), (88, 44, 133), (80, 37, 118), (74, 31, 109), (68, 27, 100), (66, 25, 93), (63, 23, 88), (61, 22, 82), (60, 21, 78), (59, 21, 74), (57, 19, 69), (56, 19, 64), (55, 18, 62), (55, 17, 59), (55, 16, 54), (55, 14, 50), (54, 13, 49), (54, 11, 48), (54, 8, 44), (54, 5, 39), (56, 3, 36), (61, 1, 33), (65, 0, 29), (59, 0, 16), (120, 57, 89), (197, 160, 201), (192, 165, 212), (190, 162, 211), (189, 163, 212), (187, 164, 213), (189, 167, 215), (189, 168, 215), (189, 168, 215), (191, 170, 217), (192, 170, 221), (190, 168, 222), (190, 168, 221), (191, 167, 220), (193, 168, 222), (193, 168, 223), (194, 168, 224), (195, 169, 226), (197, 170, 227), (198, 172, 228), (198, 173, 227), (200, 176, 229), (203, 178, 230), (205, 181, 231), (208, 185, 231), (212, 190, 232), (215, 197, 234), (221, 201, 235), (223, 203, 237), (226, 205, 238), (225, 204, 235), (223, 207, 244), (226, 195, 231), (158, 59, 68), (127, 0, 0), (143, 0, 4), (141, 0, 2), (139, 0, 0), (138, 1, 1), (137, 2, 2), (136, 1, 1), (135, 1, 0), (133, 0, 1), (130, 0, 0), (127, 0, 0), (126, 0, 0), (126, 0, 0), (126, 1, 3), (125, 2, 4), (115, 0, 1), (140, 4, 3), (207, 5, 1), (214, 0, 1), (199, 0, 0), (222, 52, 43), (255, 101, 86), (254, 96, 79), (11, 163, 226), (11, 165, 227), (13, 166, 230), (18, 166, 231), (22, 165, 231), (28, 166, 230), (29, 167, 228), (28, 165, 226), (27, 164, 228), (22, 160, 227), (12, 155, 222), (4, 149, 218), (0, 143, 213), (3, 133, 203), (2, 90, 171), (1, 60, 151), (1, 56, 146), (0, 53, 140), (1, 51, 135), (1, 50, 133), (1, 49, 133), (0, 47, 134), (1, 47, 136), (2, 46, 138), (2, 46, 138), (1, 45, 138), (2, 44, 140), (2, 46, 140), (2, 49, 139), (0, 51, 139), (0, 53, 141), (1, 52, 142), (2, 47, 129), (5, 44, 114), (7, 128, 157), (0, 154, 177), (0, 137, 168), (0, 128, 160), (0, 127, 159), (0, 125, 162), (0, 123, 162), (0, 124, 162), (0, 132, 166), (0, 132, 168), (5, 115, 160), (0, 56, 117), (138, 152, 196), (209, 179, 218), (171, 118, 192), (156, 103, 183), (155, 99, 184), (158, 99, 186), (158, 100, 189), (160, 102, 192), (164, 104, 196), (166, 107, 200), (170, 109, 199), (172, 110, 198), (173, 112, 199), (173, 110, 199), (180, 117, 203), (116, 66, 149), (87, 50, 140), (150, 112, 208), (176, 139, 231), (180, 142, 236), (180, 138, 233), (176, 129, 223), (152, 103, 194), (87, 42, 119), (39, 0, 62), (41, 0, 66), (38, 2, 62), (36, 0, 57), (51, 11, 77), (143, 100, 191), (134, 91, 194), (112, 68, 171), (98, 55, 154), (89, 45, 142), (81, 38, 125), (73, 33, 112), (67, 29, 105), (64, 27, 98), (62, 24, 92), (59, 22, 87), (57, 20, 84), (56, 21, 80), (56, 20, 76), (57, 19, 73), (55, 19, 68), (54, 19, 66), (55, 19, 65), (54, 19, 58), (53, 17, 56), (53, 15, 54), (51, 13, 50), (52, 10, 47), (53, 8, 43), (55, 6, 40), (59, 3, 38), (50, 0, 25), (85, 35, 70), (184, 149, 196), (184, 158, 207), (182, 159, 204), (184, 160, 207), (184, 160, 209), (184, 161, 211), (186, 161, 213), (185, 163, 213), (185, 163, 212), (186, 163, 213), (185, 161, 216), (184, 159, 217), (184, 160, 218), (187, 161, 218), (189, 161, 219), (189, 161, 220), (189, 160, 221), (190, 161, 222), (192, 164, 224), (194, 166, 226), (194, 166, 226), (196, 169, 226), (199, 172, 226), (202, 174, 226), (205, 178, 227), (208, 182, 228), (212, 190, 231), (217, 196, 232), (221, 201, 235), (223, 203, 237), (223, 202, 235), (220, 198, 233), (222, 202, 240), (223, 183, 213), (146, 34, 46), (137, 0, 0), (141, 1, 1), (139, 0, 0), (139, 1, 0), (139, 0, 1), (136, 0, 0), (130, 0, 0), (134, 0, 0), (144, 5, 4), (152, 11, 11), (151, 13, 11), (141, 9, 8), (128, 1, 2), (117, 0, 0), (108, 0, 0), (125, 4, 1), (205, 6, 2), (206, 0, 0), (223, 41, 37), (255, 93, 79), (247, 82, 65), (243, 71, 50), (0, 152, 218), (0, 155, 220), (0, 155, 221), (1, 156, 222), (1, 157, 223), (1, 155, 223), (2, 153, 222), (0, 151, 221), (0, 150, 219), (0, 147, 216), (0, 143, 210), (1, 137, 206), (3, 127, 202), (3, 122, 191), (3, 98, 171), (2, 64, 148), (3, 58, 142), (1, 55, 137), (0, 53, 133), (0, 52, 132), (1, 50, 132), (1, 48, 133), (2, 47, 134), (2, 46, 134), (2, 46, 135), (1, 46, 136), (1, 47, 139), (2, 47, 140), (3, 50, 141), (2, 51, 138), (2, 51, 137), (1, 49, 135), (1, 38, 112), (7, 49, 105), (3, 121, 145), (0, 116, 146), (28, 125, 157), (93, 161, 183), (144, 189, 213), (151, 195, 219), (140, 188, 214), (93, 159, 187), (28, 128, 156), (0, 110, 149), (0, 102, 152), (102, 143, 186), (253, 219, 255), (182, 136, 196), (149, 94, 172), (143, 85, 166), (141, 78, 164), (143, 77, 168), (146, 79, 175), (148, 82, 178), (152, 85, 181), (156, 89, 185), (159, 92, 188), (162, 93, 190), (163, 95, 193), (160, 90, 188), (150, 82, 176), (159, 111, 200), (173, 137, 232), (157, 117, 229), (136, 98, 214), (128, 89, 206), (128, 84, 205), (135, 86, 206), (155, 102, 218), (170, 115, 221), (99, 51, 132), (31, 0, 55), (34, 2, 57), (29, 0, 49), (80, 41, 113), (146, 102, 205), (118, 74, 181), (102, 59, 161), (92, 49, 148), (84, 41, 135), (74, 33, 118), (67, 29, 108), (64, 27, 102), (62, 25, 97), (58, 22, 91), (57, 21, 87), (56, 21, 85), (57, 21, 82), (58, 21, 78), (57, 20, 77), (55, 20, 73), (54, 20, 70), (54, 20, 68), (53, 20, 62), (53, 18, 59), (53, 17, 59), (52, 15, 55), (53, 12, 51), (53, 10, 47), (55, 9, 45), (54, 1, 40), (58, 9, 47), (164, 124, 163), (190, 160, 206), (179, 151, 200), (179, 154, 202), (179, 156, 204), (179, 157, 206), (181, 157, 209), (182, 157, 211), (181, 156, 211), (178, 155, 208), (178, 154, 208), (178, 154, 211), (179, 153, 212), (179, 151, 212), (182, 152, 214), (182, 153, 214), (183, 152, 216), (185, 152, 216), (186, 155, 216), (188, 156, 219), (190, 158, 221), (191, 159, 220), (192, 162, 219), (194, 165, 220), (198, 168, 222), (201, 171, 223), (203, 175, 224), (208, 182, 227), (212, 187, 228), (215, 193, 231), (220, 198, 234), (221, 198, 233), (222, 195, 230), (220, 194, 228), (224, 200, 243), (207, 145, 176), (130, 11, 19), (132, 0, 0), (131, 0, 0), (131, 0, 0), (129, 0, 0), (141, 0, 0), (178, 31, 29), (213, 60, 56), (238, 79, 70), (247, 90, 76), (247, 92, 76), (243, 85, 71), (225, 70, 56), (189, 45, 38), (138, 13, 13), (110, 0, 0), (183, 0, 3), (213, 21, 21), (248, 80, 74), (240, 69, 52), (234, 60, 38), (232, 55, 28), (0, 147, 214), (1, 147, 217), (0, 148, 216), (0, 148, 217), (0, 148, 217), (0, 145, 214), (0, 143, 213), (1, 140, 212), (1, 135, 209), (2, 132, 204), (2, 127, 199), (1, 122, 194), (1, 115, 187), (0, 108, 174), (0, 95, 160), (2, 70, 143), (3, 61, 141), (0, 57, 136), (1, 57, 133), (0, 54, 131), (0, 52, 132), (2, 51, 133), (2, 49, 135), (2, 48, 135), (1, 49, 135), (0, 49, 135), (1, 50, 137), (2, 49, 139), (3, 50, 138), (4, 51, 135), (3, 49, 133), (0, 45, 120), (0, 28, 86), (0, 45, 82), (9, 101, 121), (117, 163, 187), (217, 221, 244), (248, 231, 255), (249, 228, 255), (247, 228, 255), (248, 230, 255), (248, 231, 255), (222, 220, 244), (118, 161, 193), (43, 116, 154), (218, 198, 243), (233, 188, 254), (166, 115, 188), (137, 78, 155), (133, 72, 153), (130, 65, 151), (133, 64, 155), (136, 67, 161), (139, 69, 164), (144, 71, 169), (147, 74, 172), (150, 77, 177), (153, 80, 181), (153, 79, 182), (139, 62, 165), (146, 81, 186), (162, 118, 228), (125, 86, 198), (110, 66, 189), (98, 57, 180), (94, 51, 177), (96, 48, 176), (101, 50, 176), (107, 53, 178), (123, 64, 190), (145, 89, 201), (68, 30, 102), (29, 0, 45), (26, 0, 44), (102, 62, 144), (134, 88, 195), (105, 58, 166), (90, 46, 146), (83, 40, 136), (76, 34, 124), (68, 29, 112), (62, 26, 104), (60, 24, 97), (57, 22, 93), (56, 22, 90), (55, 21, 86), (56, 22, 84), (58, 22, 83), (57, 22, 82), (56, 20, 80), (56, 21, 77), (56, 20, 74), (54, 19, 71), (54, 19, 67), (53, 17, 63), (53, 17, 61), (52, 15, 58), (53, 14, 55), (52, 12, 51), (54, 11, 50), (46, 0, 40), (121, 76, 121), (189, 156, 200), (179, 149, 196), (181, 153, 202), (179, 152, 203), (177, 152, 202), (176, 152, 204), (177, 152, 206), (174, 149, 205), (173, 148, 204), (173, 148, 203), (172, 148, 205), (172, 148, 206), (172, 145, 205), (174, 142, 206), (175, 142, 207), (175, 142, 208), (176, 142, 208), (178, 143, 208), (180, 146, 210), (180, 147, 212), (183, 148, 213), (185, 151, 213), (185, 153, 212), (189, 156, 214), (192, 159, 218), (195, 163, 219), (198, 166, 219), (202, 171, 222), (205, 177, 223), (210, 183, 227), (215, 190, 231), (219, 193, 230), (218, 192, 231), (216, 192, 235), (212, 188, 232), (224, 184, 226), (183, 89, 105), (154, 24, 21), (174, 42, 37), (181, 51, 49), (185, 55, 53), (224, 89, 84), (251, 109, 100), (252, 104, 93), (247, 95, 82), (244, 86, 70), (248, 82, 65), (254, 84, 65), (255, 87, 69), (255, 89, 71), (246, 78, 66), (192, 41, 34), (160, 6, 5), (228, 55, 44), (243, 66, 44), (235, 49, 16), (232, 40, 7), (226, 32, 4), (0, 138, 206), (1, 140, 209), (1, 140, 210), (0, 140, 210), (0, 140, 210), (0, 137, 208), (0, 135, 206), (0, 132, 203), (2, 128, 199), (2, 124, 196), (2, 119, 189), (2, 111, 182), (0, 105, 171), (0, 97, 152), (0, 84, 132), (0, 65, 111), (3, 67, 131), (1, 63, 137), (0, 62, 133), (0, 60, 131), (0, 56, 132), (1, 55, 133), (1, 53, 135), (0, 52, 136), (0, 54, 135), (0, 53, 135), (2, 53, 135), (3, 53, 134), (2, 53, 133), (2, 50, 132), (1, 45, 126), (1, 38, 102), (0, 19, 64), (6, 33, 73), (151, 176, 202), (246, 226, 255), (231, 203, 245), (218, 192, 240), (216, 191, 240), (218, 192, 240), (219, 195, 237), (223, 198, 241), (233, 205, 248), (245, 219, 255), (214, 201, 239), (225, 178, 244), (218, 162, 247), (169, 110, 190), (128, 68, 145), (126, 62, 142), (126, 57, 142), (127, 57, 144), (129, 57, 147), (132, 58, 152), (137, 61, 158), (140, 62, 163), (140, 66, 166), (142, 67, 168), (137, 60, 162), (111, 42, 143), (125, 80, 191), (103, 66, 183), (87, 47, 164), (82, 40, 157), (78, 36, 152), (77, 33, 153), (77, 32, 155), (81, 32, 155), (85, 33, 155), (90, 36, 159), (114, 57, 175), (104, 52, 141), (32, 0, 43), (54, 16, 75), (127, 84, 177), (142, 96, 197), (130, 82, 181), (112, 65, 167), (88, 43, 142), (66, 25, 114), (61, 26, 102), (57, 24, 97), (54, 21, 91), (53, 21, 89), (53, 22, 89), (53, 21, 85), (54, 21, 83), (54, 22, 83), (52, 22, 82), (54, 21, 80), (53, 21, 78), (55, 21, 77), (55, 20, 75), (55, 19, 71), (52, 18, 68), (52, 18, 64), (52, 16, 60), (52, 16, 59), (52, 15, 55), (50, 8, 49), (68, 24, 68), (170, 132, 178), (178, 147, 195), (174, 147, 196), (174, 148, 199), (173, 147, 198), (173, 146, 199), (172, 146, 201), (169, 144, 200), (168, 142, 199), (169, 144, 201), (168, 144, 200), (167, 140, 197), (166, 138, 198), (166, 135, 199), (167, 133, 200), (168, 133, 201), (170, 133, 202), (171, 134, 201), (172, 135, 202), (174, 137, 205), (175, 138, 207), (178, 140, 207), (179, 142, 209), (182, 144, 210), (184, 147, 210), (187, 151, 213), (190, 155, 213), (193, 158, 214), (195, 162, 217), (200, 167, 217), (205, 173, 222), (207, 178, 228), (207, 182, 223), (215, 179, 211), (229, 165, 195), (234, 153, 167), (234, 144, 147), (247, 140, 130), (254, 140, 125), (255, 152, 138), (255, 157, 141), (255, 159, 144), (255, 159, 146), (253, 158, 146), (254, 158, 144), (251, 151, 138), (247, 144, 129), (247, 130, 116), (242, 115, 99), (238, 92, 77), (241, 74, 56), (247, 71, 53), (255, 73, 59), (226, 56, 40), (233, 60, 40), (234, 35, 11), (231, 19, 1), (224, 13, 0), (219, 5, 0), (0, 133, 200), (1, 135, 204), (3, 136, 206), (2, 136, 206), (1, 135, 206), (0, 132, 203), (1, 130, 201), (1, 127, 198), (0, 122, 192), (0, 118, 187), (0, 112, 180), (1, 105, 171), (0, 98, 163), (1, 90, 146), (3, 76, 121), (7, 74, 105), (2, 69, 109), (3, 73, 129), (1, 69, 139), (1, 65, 136), (3, 62, 135), (2, 62, 135), (2, 59, 136), (0, 56, 137), (0, 56, 137), (1, 56, 138), (2, 54, 136), (1, 53, 132), (1, 52, 130), (2, 41, 114), (5, 28, 89), (5, 26, 80), (0, 19, 61), (111, 120, 162), (230, 207, 252), (208, 173, 233), (199, 166, 231), (199, 160, 231), (203, 160, 232), (205, 162, 232), (206, 163, 234), (210, 168, 235), (212, 175, 236), (219, 186, 242), (227, 186, 253), (213, 150, 248), (215, 142, 254), (190, 119, 221), (131, 67, 145), (126, 60, 139), (126, 55, 141), (127, 54, 141), (125, 52, 140), (125, 50, 144), (128, 48, 148), (130, 50, 150), (128, 52, 151), (125, 50, 148), (112, 35, 133), (91, 28, 125), (96, 55, 159), (72, 36, 139), (68, 30, 131), (64, 26, 128), (63, 23, 127), (65, 23, 130), (66, 23, 132), (67, 22, 134), (71, 22, 138), (77, 25, 140), (87, 31, 141), (99, 45, 144), (116, 72, 158), (139, 97, 193), (134, 90, 204), (132, 85, 197), (135, 85, 194), (137, 86, 194), (129, 77, 183), (101, 56, 152), (60, 28, 103), (49, 19, 88), (51, 20, 88), (50, 20, 86), (50, 21, 85), (48, 19, 83), (49, 20, 81), (50, 19, 80), (50, 19, 80), (52, 19, 78), (53, 19, 77), (54, 19, 77), (54, 19, 76), (54, 19, 75), (54, 19, 72), (53, 18, 68), (52, 18, 64), (52, 16, 62), (52, 16, 58), (43, 4, 47), (116, 77, 123), (182, 149, 196), (171, 141, 191), (171, 144, 196), (170, 143, 195), (167, 140, 193), (166, 139, 194), (165, 138, 194), (164, 138, 194), (163, 138, 195), (161, 136, 194), (160, 135, 193), (158, 131, 191), (160, 129, 193), (160, 127, 193), (158, 124, 192), (160, 123, 192), (161, 122, 192), (163, 123, 193), (165, 124, 194), (168, 126, 197), (171, 128, 200), (172, 130, 200), (174, 132, 199), (177, 134, 201), (178, 138, 204), (180, 141, 204), (184, 143, 205), (189, 145, 208), (191, 147, 210), (190, 151, 210), (190, 155, 209), (205, 156, 194), (226, 151, 166), (239, 143, 142), (252, 139, 125), (255, 143, 124), (255, 145, 128), (255, 151, 133), (255, 153, 140), (255, 154, 141), (253, 154, 138), (253, 154, 140), (251, 156, 144), (250, 157, 147), (252, 158, 150), (255, 164, 155), (254, 167, 155), (253, 166, 153), (254, 167, 155), (251, 162, 145), (243, 140, 123), (239, 100, 91), (241, 66, 55), (243, 55, 33), (230, 35, 15), (224, 7, 0), (221, 0, 0), (220, 0, 0), (216, 0, 1), (0, 130, 196), (1, 131, 198), (3, 132, 198), (1, 130, 197), (0, 128, 196), (0, 126, 194), (2, 124, 194), (2, 122, 190), (2, 117, 180), (0, 109, 172), (0, 103, 166), (1, 100, 160), (0, 96, 155), (2, 86, 139), (4, 78, 119), (9, 100, 127), (2, 64, 88), (3, 64, 91), (8, 71, 120), (8, 73, 143), (3, 73, 140), (0, 68, 134), (1, 65, 135), (1, 62, 137), (0, 60, 135), (2, 58, 133), (1, 55, 130), (1, 50, 119), (1, 39, 104), (4, 48, 103), (7, 86, 122), (4, 115, 141), (34, 121, 158), (192, 182, 234), (192, 153, 224), (179, 130, 216), (177, 132, 214), (172, 129, 215), (174, 127, 217), (177, 127, 221), (184, 129, 227), (191, 138, 231), (192, 145, 230), (197, 153, 237), (210, 156, 252), (206, 131, 250), (207, 122, 254), (208, 126, 251), (154, 83, 175), (125, 57, 137), (126, 56, 139), (124, 52, 138), (121, 48, 136), (118, 42, 134), (117, 38, 132), (116, 34, 131), (111, 31, 130), (105, 29, 125), (85, 10, 99), (74, 18, 107), (71, 34, 127), (57, 24, 107), (54, 21, 101), (52, 17, 100), (52, 15, 102), (54, 14, 107), (55, 14, 113), (58, 14, 117), (63, 16, 122), (68, 19, 125), (76, 21, 126), (91, 38, 142), (129, 83, 203), (109, 67, 195), (97, 53, 184), (94, 45, 178), (94, 41, 171), (94, 39, 161), (96, 39, 158), (105, 50, 167), (102, 50, 150), (56, 20, 96), (40, 17, 77), (44, 19, 78), (45, 18, 78), (45, 17, 75), (46, 17, 76), (47, 17, 76), (47, 17, 74), (50, 17, 76), (48, 17, 76), (48, 18, 75), (51, 19, 75), (53, 20, 73), (52, 19, 73), (52, 19, 70), (52, 20, 67), (52, 18, 65), (50, 14, 59), (53, 17, 62), (155, 119, 167), (174, 145, 193), (168, 141, 189), (167, 140, 190), (164, 138, 191), (161, 133, 189), (159, 132, 189), (159, 131, 187), (159, 131, 187), (154, 128, 186), (152, 126, 185), (150, 122, 183), (150, 120, 182), (152, 119, 183), (151, 117, 183), (152, 115, 185), (154, 114, 185), (156, 114, 185), (157, 113, 185), (158, 114, 186), (161, 117, 189), (165, 118, 191), (166, 119, 192), (168, 121, 192), (171, 122, 192), (172, 123, 193), (174, 125, 193), (177, 127, 194), (181, 130, 198), (179, 131, 199), (189, 135, 179), (220, 136, 153), (242, 138, 131), (255, 135, 115), (255, 137, 121), (255, 142, 122), (254, 145, 128), (254, 148, 133), (254, 149, 134), (253, 149, 132), (253, 148, 132), (251, 149, 133), (253, 152, 137), (254, 153, 141), (252, 158, 146), (254, 161, 151), (253, 157, 146), (253, 155, 142), (254, 157, 143), (253, 163, 149), (254, 167, 151), (255, 167, 157), (253, 166, 157), (246, 148, 135), (238, 85, 72), (214, 6, 2), (224, 0, 0), (221, 1, 2), (217, 1, 1), (213, 1, 2), (0, 128, 192), (0, 128, 192), (2, 128, 192), (1, 125, 190), (0, 123, 189), (1, 122, 187), (0, 119, 184), (0, 116, 181), (2, 111, 172), (0, 103, 163), (0, 99, 155), (2, 97, 150), (1, 94, 148), (0, 84, 127), (5, 86, 115), (6, 84, 114), (2, 50, 74), (2, 44, 56), (2, 43, 61), (4, 52, 79), (4, 65, 105), (4, 73, 125), (3, 71, 128), (4, 67, 127), (3, 66, 122), (1, 62, 115), (1, 57, 105), (1, 55, 91), (8, 70, 108), (9, 120, 155), (4, 148, 178), (0, 152, 179), (81, 161, 205), (190, 148, 219), (177, 136, 203), (206, 172, 224), (223, 191, 236), (222, 195, 239), (221, 194, 239), (215, 183, 235), (196, 153, 220), (174, 117, 212), (171, 110, 222), (176, 114, 226), (198, 129, 241), (199, 114, 246), (200, 108, 248), (203, 113, 250), (195, 110, 236), (139, 67, 162), (121, 54, 135), (119, 48, 134), (113, 42, 127), (101, 29, 113), (89, 16, 102), (79, 8, 96), (75, 5, 95), (70, 3, 88), (59, 1, 68), (54, 8, 81), (53, 19, 92), (45, 16, 87), (43, 11, 88), (44, 8, 89), (45, 7, 92), (47, 6, 96), (49, 6, 104), (53, 8, 110), (59, 11, 117), (64, 15, 121), (71, 18, 122), (74, 24, 126), (76, 29, 154), (78, 33, 170), (75, 30, 166), (73, 22, 164), (72, 14, 163), (71, 10, 157), (68, 7, 150), (71, 5, 142), (89, 19, 144), (87, 26, 132), (46, 15, 76), (38, 19, 70), (42, 18, 73), (43, 18, 73), (44, 16, 74), (45, 16, 74), (45, 16, 73), (47, 16, 74), (46, 17, 73), (46, 17, 72), (47, 16, 71), (48, 16, 69), (48, 17, 69), (48, 18, 68), (49, 18, 67), (51, 17, 65), (43, 10, 57), (82, 48, 96), (172, 139, 190), (165, 137, 188), (163, 135, 186), (161, 133, 184), (158, 129, 183), (154, 125, 182), (153, 124, 182), (152, 122, 180), (150, 120, 177), (145, 118, 175), (143, 115, 174), (142, 111, 174), (142, 109, 174), (142, 106, 173), (143, 105, 174), (145, 104, 175), (146, 103, 175), (147, 103, 175), (148, 102, 175), (150, 103, 176), (153, 105, 178), (154, 105, 178), (157, 105, 179), (159, 105, 179), (160, 105, 178), (163, 106, 178), (163, 107, 180), (163, 108, 179), (169, 106, 175), (204, 119, 155), (241, 130, 121), (255, 130, 113), (255, 132, 114), (255, 136, 120), (254, 137, 120), (253, 137, 120), (252, 140, 123), (253, 141, 125), (252, 136, 121), (254, 141, 125), (253, 144, 128), (252, 146, 131), (252, 147, 133), (255, 151, 138), (254, 154, 140), (252, 153, 140), (253, 152, 138), (253, 152, 138), (254, 153, 139), (253, 154, 140), (251, 152, 139), (251, 152, 136), (252, 153, 137), (254, 159, 144), (255, 162, 148), (241, 126, 111), (219, 34, 36), (220, 0, 2), (216, 2, 3), (210, 1, 1)
);

end package pmod_lcd_pkg;
-------------------------------------------------------------------------------
package body pmod_lcd_pkg is

end package body pmod_lcd_pkg;